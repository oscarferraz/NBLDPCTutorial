`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.01.2020 18:13:04
// Design Name: 
// Module Name: test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test();
reg clk,reset;
reg [5:0]in;
wire[5:0]out;
wire out_enable;
integer handle1;
minmaxdecoding rgr(clk,reset,in,out,out_enable);

initial
begin

 handle1 = $fopen("file1.out");

end

always@(posedge clk) begin
$fdisplay(handle1,"%d",out);
end

initial begin
#13000000 $finish;
end


initial
clk=1'b0;
initial
reset=0;

initial
#110 reset=1;
initial
#120 reset=0;

initial
begin
 #100 in=6'd2;
#470 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd2;

#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd18;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd18;
#400 in=6'd18;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd17;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd15;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd12;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd13;
#400 in=6'd6;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd13;
#400 in=6'd6;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd17;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd12;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd18;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd13;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd19;
#400 in=6'd13;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd7;
#400 in=6'd15;
#400 in=6'd14;
#400 in=6'd21;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd16;
#400 in=6'd23;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd18;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd12;
#400 in=6'd19;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd18;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd19;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd18;
#400 in=6'd17;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd11;
#400 in=6'd18;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd11;
#400 in=6'd18;
#400 in=6'd15;
#400 in=6'd22;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd16;
#400 in=6'd17;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd16;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd17;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd17;
#400 in=6'd3;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd15;
#400 in=6'd8;
#400 in=6'd18;
#400 in=6'd10;
#400 in=6'd20;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd11;
#400 in=6'd19;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd19;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd13;
#400 in=6'd4;
#400 in=6'd14;
#400 in=6'd7;
#400 in=6'd16;
#400 in=6'd7;
#400 in=6'd16;
#400 in=6'd9;
#400 in=6'd18;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd12;
#400 in=6'd18;
#400 in=6'd16;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd19;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd19;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd16;
#400 in=6'd23;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd18;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd17;
#400 in=6'd15;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd17;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd12;
#400 in=6'd20;
#400 in=6'd14;
#400 in=6'd22;
#400 in=6'd17;
#400 in=6'd25;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd18;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd18;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd17;
#400 in=6'd8;
#400 in=6'd19;
#400 in=6'd1;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd19;
#400 in=6'd9;
#400 in=6'd20;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd17;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd17;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd18;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd16;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd14;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd14;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd1;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd17;
#400 in=6'd22;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd16;
#400 in=6'd22;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd17;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd17;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd18;
#400 in=6'd6;
#400 in=6'd15;
#400 in=6'd12;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd16;
#400 in=6'd23;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd14;
#400 in=6'd19;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd14;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd15;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd18;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd20;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd17;
#400 in=6'd17;
#400 in=6'd19;
#400 in=6'd23;
#400 in=6'd25;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd17;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd19;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd22;
#400 in=6'd2;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd16;
#400 in=6'd5;
#400 in=6'd14;
#400 in=6'd6;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd14;
#400 in=6'd11;
#400 in=6'd20;
#400 in=6'd9;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd14;
#400 in=6'd19;
#400 in=6'd16;
#400 in=6'd20;
#400 in=6'd18;
#400 in=6'd23;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd20;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd15;
#400 in=6'd20;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd17;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd16;
#400 in=6'd16;
#400 in=6'd18;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd15;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd17;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd18;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd17;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd18;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd14;
#400 in=6'd1;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd15;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd1;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd17;
#400 in=6'd18;
#400 in=6'd21;
#400 in=6'd23;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd22;
#400 in=6'd16;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd13;
#400 in=6'd20;
#400 in=6'd1;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd12;
#400 in=6'd20;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd12;
#400 in=6'd19;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd15;
#400 in=6'd10;
#400 in=6'd19;
#400 in=6'd6;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd18;
#400 in=6'd12;
#400 in=6'd21;
#400 in=6'd16;
#400 in=6'd24;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd13;
#400 in=6'd19;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd18;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd19;
#400 in=6'd12;
#400 in=6'd18;
#400 in=6'd18;
#400 in=6'd25;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd18;
#400 in=6'd7;
#400 in=6'd15;
#400 in=6'd14;
#400 in=6'd21;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd18;
#400 in=6'd20;
#400 in=6'd22;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd17;
#400 in=6'd24;
#400 in=6'd18;
#400 in=6'd24;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd13;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd15;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd12;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd17;
#400 in=6'd16;
#400 in=6'd20;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd13;
#400 in=6'd18;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd13;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd17;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd16;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd19;
#400 in=6'd18;
#400 in=6'd22;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd15;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd18;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd15;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd14;
#400 in=6'd20;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd14;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd16;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd19;
#400 in=6'd21;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd15;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd15;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd20;
#400 in=6'd11;
#400 in=6'd14;
#400 in=6'd20;
#400 in=6'd23;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd5;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd1;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd11;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd7;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd12;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd9;
#400 in=6'd16;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd13;
#400 in=6'd15;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd8;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd13;
#400 in=6'd16;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd1;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd9;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd10;
#400 in=6'd4;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd7;
#400 in=6'd15;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd2;
#400 in=6'd10;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd16;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd11;
#400 in=6'd17;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd14;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd10;
#400 in=6'd12;
#400 in=6'd0;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd5;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd19;
#400 in=6'd7;
#400 in=6'd14;
#400 in=6'd13;
#400 in=6'd21;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd5;
#400 in=6'd1;
#400 in=6'd6;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd4;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd13;
#400 in=6'd8;
#400 in=6'd13;
#400 in=6'd11;
#400 in=6'd16;
#400 in=6'd12;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd6;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd9;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd9;
#400 in=6'd15;
#400 in=6'd2;
#400 in=6'd5;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd8;
#400 in=6'd10;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd8;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd1;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd6;
#400 in=6'd12;
#400 in=6'd2;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd7;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd11;
#400 in=6'd10;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd16;
#400 in=6'd15;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd19;
#400 in=6'd17;
#400 in=6'd0;
#400 in=6'd2;
#400 in=6'd7;
#400 in=6'd9;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd9;
#400 in=6'd11;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd11;
#400 in=6'd13;
#400 in=6'd0;
#400 in=6'd1;
#400 in=6'd1;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd5;
#400 in=6'd5;
#400 in=6'd6;
#400 in=6'd2;
#400 in=6'd3;
#400 in=6'd3;
#400 in=6'd4;
#400 in=6'd6;
#400 in=6'd7;
#400 in=6'd7;
#400 in=6'd8;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd15;
#400 in=6'd19;
#400 in=6'd13;
#400 in=6'd17;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd10;
#400 in=6'd14;
#400 in=6'd2;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd14;
#400 in=6'd18;
#400 in=6'd12;
#400 in=6'd16;
#400 in=6'd5;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd17;
#400 in=6'd21;
#400 in=6'd15;
#400 in=6'd19;
#400 in=6'd0;
#400 in=6'd9;
#400 in=6'd3;
#400 in=6'd12;
#400 in=6'd4;
#400 in=6'd13;
#400 in=6'd7;
#400 in=6'd16;
#400 in=6'd6;
#400 in=6'd15;
#400 in=6'd9;
#400 in=6'd18;
#400 in=6'd10;
#400 in=6'd19;
#400 in=6'd13;
#400 in=6'd22;
#400 in=6'd0;
#400 in=6'd7;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd3;
#400 in=6'd10;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd5;
#400 in=6'd12;
#400 in=6'd10;
#400 in=6'd17;
#400 in=6'd8;
#400 in=6'd15;
#400 in=6'd13;
#400 in=6'd20;
#400 in=6'd0;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd3;
#400 in=6'd7;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd3;
#400 in=6'd8;
#400 in=6'd6;
#400 in=6'd10;
#400 in=6'd7;
#400 in=6'd11;
#400 in=6'd9;
#400 in=6'd13;
#400 in=6'd1;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd2;
#400 in=6'd4;
#400 in=6'd3;
#400 in=6'd6;
#400 in=6'd0;
#400 in=6'd3;
#400 in=6'd2;
#400 in=6'd5;

end
initial
begin
forever 
#200 clk=~clk;
end
endmodule
//create_clock -period 12.000 -name clk -waveform {0.000 6.000} -add [get_ports clk]
//create_clock -period 12.000 -name clk -waveform {0.000 6.000} -add [get_ports clk]
