
module minmaxdecoding(gamma,reset,clk,beta);
parameter Gammalen=5;
parameter addrlen=2;
parameter collen=9;
parameter rowlen=8;
parameter Nbits=3;
parameter QQ=7;
input[Gammalen-1:0]gamma;
input reset;
input clk;
output reg[Gammalen:0] beta;
reg[10:0]address_index,address_index1,address_index2;

/* ALL FUNCTIONS ARE DEFINED BELOW*/

function[Gammalen:0] max;
    input[Gammalen:0] p,q;
    if(p<q) max=q;
    else max=p;
    endfunction
    
function[Gammalen:0] min;
        input[Gammalen:0] p,q;
        if(p<q) min=p;
        else min=q;
        endfunction  


/* ALL THE TASKS ARE DEFINED BELOW*/



task mul_gf;// this one defines the multiplication for gf(4)  
input[2:0] A;
input[2:0]B;
output [2:0]Y;
begin

	
Y={(A[2]&B[2])^(A[2]&B[0])^(A[1]&B[1])^(A[0]&B[2]),(A[2]&B[2])^(A[2]&B[1])^(A[1]&B[2])^(A[1]&B[0])^(A[0]&B[1]),(A[2]&B[1])^(A[1]&B[2])^(A[0]&B[0])};

end
endtask

task add_gf;// this one defines the addition for gf(4)   
input[2:0] A;//this is simply xor operation of bits
input [2:0]Be;
output[2:0] out;
begin
out[0]=A[0]^Be[0];
out[1]=A[1]^Be[1];
out[2]=A[2]^Be[2];
end
endtask


task inv_gf;// this task computes the multiplicative inverse of a given number
input[2:0] A;
output [2:0]  out;
begin
//out= expq[(7 - logq[A])];
//if(A == 0) out=0;
//	if(A == 1) out=1;
	
if(A==3'd0)
out=3'd0;
else if(A==3'd1)
out=3'd1;
else if(A<3'd5)
out=A+3'd3;
else
out=A-3'd3;
end
endtask





/* ALL DEFINED CONSTANTS ARE BELOW*/
`define gammaIn 6'd0
`define alpha_Init 6'd1
`define processing_state 6'd2
`define F_init1 6'd3
`define processing_state1 6'd4
`define B_init1 6'd5
`define processing_state2 6'd6
`define processing_state3 6'd7
`define Alphadecide 6'd8
`define F_init2 6'd9
`define processing_state4 6'd10
`define processing_state5 6'd11
`define Alphadecide1 6'd12
`define B_init2 6'd13
`define s39 6'd14
`define BETA1 6'd15
`define BETA2 6'd16
`define BETA3 6'd17
`define BETAOUT 6'd18 
`define processing_state7 6'd19
`define processing_state6 6'd20
`define WAIT 6'd21
`define F_init21 6'd22
`define B_init21 6'd23
`define BETA31 6'd24
`define processing_state8 6'd25
`define FindMin 6'd26
`define FixAlpha 6'd27
`define GammaFix 6'd28
`define processing_statex 6'd29
`define temporary_state_1 6'd30
`define BETADECIDE 6'd31
`define temporary_state_2 6'd32
`define BETAOUT1 6'd33
`define BETAOUT2 6'd34
`define s1 6'd40
`define s2 6'd41
`define s3 6'd42
`define s4 6'd43
`define s5 6'd44
`define s6 6'd45
`define s7 6'd46
`define ITERATION 4'd10

/* ALL REGISTER DECLARATIONS ARE BELOW FOR CHECK NODE PROCESSING*/
reg[5:0]state;
//reg weA,weB;
reg[1:0] expanded_address;////////////////////////////
//reg[addrlen:0] addrAR,addrAW,addrBR,addrBW;
//reg[Gammalen:0]dinA,dinB;
//wire[Gammalen:0]doutA,doutB;
reg[rowlen:0]row,row2,reading_row;
reg[Nbits:0]H[255:0][383:0];
reg[collen:0]col,col1,col2;
reg[Gammalen:0]Gamma[QQ:0][383:0];
reg[Gammalen:0]F[QQ:0][2:0][255:0];/////BASED ON RW AND CW
reg[Gammalen:0]B[QQ:0][2:0][255:0];////// BASED ON RW AND CW
reg[Nbits:0]x,y,c,a,reading_a,inv_val,mul_val,mul_val1,s,b;
reg index_VN[255:0][383:0];
reg[collen:0]col_row[255:0][2:0];
reg[rowlen:0]row_col[1:0][383:0];
reg[Gammalen:0]AlphaSet[QQ:0][255:0];
reg[Gammalen:0]min_F[255:0][QQ:0],max_F[255:0][QQ:0];
reg[Gammalen:0]min_B[255:0][QQ:0],max_B[255:0][QQ:0],unused_variable;
reg[1:0]index_CN[255:0][383:0];
reg[1:0]temp_address;

/* ALL THE ABOVE ARE FOR CHECK NODE PROCESSING ONLY*/

/* the iter register*/
reg[3:0]iter;

/* THE BELOW ARE THE REGISTERS REQD FOR VARIABLE NODE PROCESSING*/

reg index_v,index;
reg[collen:0]betaset[QQ:0];
reg[collen:0]ALPHA_t[QQ:0];
reg [6:0]tempa[QQ:0][383:0];
reg [6:0]tempm[QQ:0][383:0];
reg [9:0]m,p,row_;
reg [Nbits:0]magic_,magicin;
reg [Nbits:0]minindex[3:0][383:0];
reg [Nbits:0]minindex_[3:0][383:0];

reg [10:0]r,t;

   reg           weA[767:0];
    reg  [addrlen:0]    addrAW[767:0];
    reg  [addrlen:0]    addrAR[767:0];
    reg  [Gammalen:0]   dinA[767:0];
    wire [Gammalen:0]   doutA[767:0];
genvar i;
    generate
    for(i=0;i<768;i=i+1)
    begin
    bram alpha(clk,weA[i],addrAW[i],addrAR[i],dinA[i],doutA[i]);
    end
    endgenerate


    reg          weB[767:0];
    reg  [addrlen:0]    addrBW[767:0];
    reg  [addrlen:0]    addrBR[767:0];
    reg  [Gammalen:0]   dinB[767:0];
    wire [Gammalen:0]   doutB[767:0];
genvar J;
    generate
    for(J=0;J<768;J=J+1)
    begin
    bram BETA(clk,weB[J],addrBW[J],addrBR[J],dinB[J],doutB[J]);
    end
    endgenerate




always@(posedge clk) begin
if(reset) begin
state=`gammaIn;
iter=`ITERATION;


//logq[0]=0;
//logq[1]=0;
//logq[2]=1;
//logq[3]=3;
//logq[4]=2;
//logq[5]=6;
//logq[6]=4;
//logq[7]=5;
//expq[0]=1;
//expq[1]=2;
//expq[2]=4;
//expq[3]=3;
//expq[4]=6;
//expq[5]=7;
//expq[6]=5;












/* BELOW IS THE INITIALIZATION FOR THE H MATRIX*/
H[0][0]=1;
H[0][1]=1;
H[0][256]=1;
H[1][1]=1;
H[1][2]=1;
H[1][257]=1;
H[2][2]=1;
H[2][3]=1;
H[2][258]=1;
H[3][3]=1;
H[3][4]=1;
H[3][259]=1;
H[4][4]=1;
H[4][5]=1;
H[4][260]=1;
H[5][5]=1;
H[5][6]=3;
H[5][261]=1;
H[6][6]=1;
H[6][7]=1;
H[6][262]=2;
H[7][7]=1;
H[7][8]=6;
H[7][263]=1;
H[8][8]=1;
H[8][9]=1;
H[8][264]=1;
H[9][9]=3;
H[9][10]=1;
H[9][265]=3;
H[10][10]=1;
H[10][11]=1;
H[10][266]=3;
H[11][11]=2;
H[11][12]=1;
H[11][267]=1;
H[12][12]=1;
H[12][13]=1;
H[12][268]=1;
H[13][13]=1;
H[13][14]=2;
H[13][269]=1;
H[14][14]=1;
H[14][15]=1;
H[14][270]=1;
H[15][15]=1;
H[15][16]=1;
H[15][271]=1;
H[16][16]=1;
H[16][17]=1;
H[16][272]=2;
H[17][17]=1;
H[17][18]=1;
H[17][273]=7;
H[18][18]=1;
H[18][19]=1;
H[18][274]=1;
H[19][19]=1;
H[19][20]=1;
H[19][275]=1;
H[20][20]=1;
H[20][21]=1;
H[20][276]=6;
H[21][21]=1;
H[21][22]=1;
H[21][277]=1;
H[22][22]=1;
H[22][23]=1;
H[22][278]=1;
H[23][23]=1;
H[23][24]=1;
H[23][279]=1;
H[24][24]=1;
H[24][25]=1;
H[24][280]=1;
H[25][25]=3;
H[25][26]=1;
H[25][281]=1;
H[26][26]=3;
H[26][27]=1;
H[26][282]=1;
H[27][27]=2;
H[27][28]=1;
H[27][283]=1;
H[28][28]=1;
H[28][29]=1;
H[28][284]=1;
H[29][29]=1;
H[29][30]=3;
H[29][285]=3;
H[30][30]=3;
H[30][31]=3;
H[30][286]=1;
H[31][31]=1;
H[31][32]=1;
H[31][287]=6;
H[32][32]=1;
H[32][33]=1;
H[32][288]=1;
H[33][33]=1;
H[33][34]=2;
H[33][289]=1;
H[34][34]=1;
H[34][35]=1;
H[34][290]=1;
H[35][35]=3;
H[35][36]=3;
H[35][291]=1;
H[36][36]=1;
H[36][37]=1;
H[36][292]=2;
H[37][37]=1;
H[37][38]=1;
H[37][293]=1;
H[38][38]=1;
H[38][39]=1;
H[38][294]=3;
H[39][39]=2;
H[39][40]=1;
H[39][295]=1;
H[40][40]=7;
H[40][41]=1;
H[40][296]=7;
H[41][41]=1;
H[41][42]=1;
H[41][297]=1;
H[42][42]=1;
H[42][43]=2;
H[42][298]=1;
H[43][43]=1;
H[43][44]=1;
H[43][299]=1;
H[44][44]=1;
H[44][45]=1;
H[44][300]=1;
H[45][45]=1;
H[45][46]=1;
H[45][301]=1;
H[46][46]=1;
H[46][47]=1;
H[46][302]=2;
H[47][47]=2;
H[47][48]=1;
H[47][303]=1;
H[48][48]=3;
H[48][49]=1;
H[48][304]=1;
H[49][49]=1;
H[49][50]=1;
H[49][305]=1;
H[50][50]=1;
H[50][51]=3;
H[50][306]=3;
H[51][51]=3;
H[51][52]=1;
H[51][307]=3;
H[52][52]=1;
H[52][53]=1;
H[52][308]=1;
H[53][53]=1;
H[53][54]=3;
H[53][309]=1;
H[54][54]=1;
H[54][55]=1;
H[54][310]=1;
H[55][55]=1;
H[55][56]=1;
H[55][311]=1;
H[56][56]=1;
H[56][57]=1;
H[56][312]=1;
H[57][57]=1;
H[57][58]=1;
H[57][313]=1;
H[58][58]=1;
H[58][59]=1;
H[58][314]=7;
H[59][59]=1;
H[59][60]=2;
H[59][315]=1;
H[60][60]=1;
H[60][61]=1;
H[60][316]=1;
H[61][61]=2;
H[61][62]=1;
H[61][317]=1;
H[62][62]=1;
H[62][63]=6;
H[62][318]=1;
H[63][63]=1;
H[63][64]=2;
H[63][319]=1;
H[64][64]=1;
H[64][65]=2;
H[64][320]=1;
H[65][65]=1;
H[65][66]=1;
H[65][321]=1;
H[66][66]=1;
H[66][67]=1;
H[66][322]=1;
H[67][67]=1;
H[67][68]=1;
H[67][323]=1;
H[68][68]=1;
H[68][69]=3;
H[68][324]=3;
H[69][69]=1;
H[69][70]=7;
H[69][325]=1;
H[70][70]=1;
H[70][71]=1;
H[70][326]=1;
H[71][71]=1;
H[71][72]=6;
H[71][327]=1;
H[72][72]=3;
H[72][73]=1;
H[72][328]=1;
H[73][73]=1;
H[73][74]=3;
H[73][329]=3;
H[74][74]=1;
H[74][75]=1;
H[74][330]=2;
H[75][75]=1;
H[75][76]=1;
H[75][331]=1;
H[76][76]=1;
H[76][77]=1;
H[76][332]=3;
H[77][77]=1;
H[77][78]=2;
H[77][333]=1;
H[78][78]=3;
H[78][79]=1;
H[78][334]=1;
H[79][79]=1;
H[79][80]=6;
H[79][335]=1;
H[80][80]=1;
H[80][81]=3;
H[80][336]=1;
H[81][81]=1;
H[81][82]=2;
H[81][337]=1;
H[82][82]=1;
H[82][83]=1;
H[82][338]=1;
H[83][83]=1;
H[83][84]=1;
H[83][339]=1;
H[84][84]=1;
H[84][85]=1;
H[84][340]=1;
H[85][85]=7;
H[85][86]=7;
H[85][341]=1;
H[86][86]=1;
H[86][87]=2;
H[86][342]=1;
H[87][87]=1;
H[87][88]=1;
H[87][343]=1;
H[88][88]=1;
H[88][89]=1;
H[88][344]=6;
H[89][89]=1;
H[89][90]=1;
H[89][345]=1;
H[90][90]=1;
H[90][91]=1;
H[90][346]=1;
H[91][91]=6;
H[91][92]=1;
H[91][347]=1;
H[92][92]=1;
H[92][93]=1;
H[92][348]=1;
H[93][93]=1;
H[93][94]=6;
H[93][349]=1;
H[94][94]=1;
H[94][95]=2;
H[94][350]=1;
H[95][95]=1;
H[95][96]=1;
H[95][351]=1;
H[96][96]=2;
H[96][97]=1;
H[96][352]=1;
H[97][97]=1;
H[97][98]=1;
H[97][353]=2;
H[98][98]=1;
H[98][99]=1;
H[98][354]=1;
H[99][99]=1;
H[99][100]=1;
H[99][355]=1;
H[100][100]=1;
H[100][101]=6;
H[100][356]=1;
H[101][101]=3;
H[101][102]=1;
H[101][357]=3;
H[102][102]=1;
H[102][103]=1;
H[102][358]=3;
H[103][103]=1;
H[103][104]=2;
H[103][359]=1;
H[104][104]=1;
H[104][105]=1;
H[104][360]=1;
H[105][105]=3;
H[105][106]=1;
H[105][361]=1;
H[106][106]=1;
H[106][107]=7;
H[106][362]=1;
H[107][107]=1;
H[107][108]=1;
H[107][363]=7;
H[108][108]=1;
H[108][109]=1;
H[108][364]=6;
H[109][109]=1;
H[109][110]=1;
H[109][365]=2;
H[110][110]=1;
H[110][111]=1;
H[110][366]=1;
H[111][111]=1;
H[111][112]=3;
H[111][367]=1;
H[112][112]=1;
H[112][113]=1;
H[112][368]=1;
H[113][113]=1;
H[113][114]=1;
H[113][369]=1;
H[114][114]=1;
H[114][115]=1;
H[114][370]=2;
H[115][115]=2;
H[115][116]=1;
H[115][371]=1;
H[116][116]=1;
H[116][117]=1;
H[116][372]=3;
H[117][117]=6;
H[117][118]=1;
H[117][373]=1;
H[118][118]=1;
H[118][119]=1;
H[118][374]=7;
H[119][119]=2;
H[119][120]=1;
H[119][375]=1;
H[120][120]=3;
H[120][121]=1;
H[120][376]=3;
H[121][121]=1;
H[121][122]=1;
H[121][377]=1;
H[122][122]=1;
H[122][123]=1;
H[122][378]=1;
H[123][123]=3;
H[123][124]=1;
H[123][379]=1;
H[124][124]=1;
H[124][125]=1;
H[124][380]=1;
H[125][125]=1;
H[125][126]=1;
H[125][381]=1;
H[126][126]=1;
H[126][127]=2;
H[126][382]=1;
H[127][0]=1;
H[127][127]=2;
H[127][383]=1;
H[128][128]=1;
H[128][129]=1;
H[128][334]=1;
H[129][129]=1;
H[129][130]=1;
H[129][268]=1;
H[130][130]=3;
H[130][131]=3;
H[130][359]=1;
H[131][131]=1;
H[131][132]=1;
H[131][342]=1;
H[132][132]=1;
H[132][133]=1;
H[132][257]=3;
H[133][133]=1;
H[133][134]=1;
H[133][320]=6;
H[134][134]=1;
H[134][135]=3;
H[134][297]=3;
H[135][135]=1;
H[135][136]=1;
H[135][264]=6;
H[136][136]=1;
H[136][137]=1;
H[136][326]=1;
H[137][137]=3;
H[137][138]=1;
H[137][355]=1;
H[138][138]=3;
H[138][139]=1;
H[138][289]=3;
H[139][139]=3;
H[139][140]=1;
H[139][314]=1;
H[140][140]=1;
H[140][141]=1;
H[140][336]=1;
H[141][141]=1;
H[141][142]=1;
H[141][256]=2;
H[142][142]=1;
H[142][143]=1;
H[142][277]=1;
H[143][143]=2;
H[143][144]=1;
H[143][350]=1;
H[144][144]=3;
H[144][145]=1;
H[144][307]=1;
H[145][145]=1;
H[145][146]=1;
H[145][266]=1;
H[146][146]=3;
H[146][147]=1;
H[146][363]=1;
H[147][147]=3;
H[147][148]=3;
H[147][300]=1;
H[148][148]=1;
H[148][149]=1;
H[148][259]=1;
H[149][149]=1;
H[149][150]=1;
H[149][325]=1;
H[150][150]=1;
H[150][151]=2;
H[150][293]=1;
H[151][151]=1;
H[151][152]=1;
H[151][367]=1;
H[152][152]=1;
H[152][153]=2;
H[152][269]=1;
H[153][153]=1;
H[153][154]=1;
H[153][278]=2;
H[154][154]=1;
H[154][155]=6;
H[154][339]=1;
H[155][155]=1;
H[155][156]=2;
H[155][322]=1;
H[156][156]=1;
H[156][157]=1;
H[156][261]=3;
H[157][157]=1;
H[157][158]=1;
H[157][356]=2;
H[158][158]=2;
H[158][159]=1;
H[158][305]=1;
H[159][159]=6;
H[159][160]=1;
H[159][272]=1;
H[160][160]=1;
H[160][161]=2;
H[160][371]=1;
H[161][161]=1;
H[161][162]=1;
H[161][344]=1;
H[162][162]=1;
H[162][163]=2;
H[162][315]=1;
H[163][163]=6;
H[163][164]=1;
H[163][294]=1;
H[164][164]=1;
H[164][165]=6;
H[164][351]=1;
H[165][165]=1;
H[165][166]=1;
H[165][262]=1;
H[166][166]=1;
H[166][167]=3;
H[166][378]=1;
H[167][167]=7;
H[167][168]=1;
H[167][288]=6;
H[168][168]=1;
H[168][169]=6;
H[168][330]=1;
H[169][169]=1;
H[169][170]=1;
H[169][343]=2;
H[170][170]=1;
H[170][171]=1;
H[170][279]=1;
H[171][171]=1;
H[171][172]=2;
H[171][374]=1;
H[172][172]=1;
H[172][173]=1;
H[172][265]=1;
H[173][173]=1;
H[173][174]=1;
H[173][337]=1;
H[174][174]=1;
H[174][175]=1;
H[174][285]=1;
H[175][175]=1;
H[175][176]=1;
H[175][302]=2;
H[176][176]=1;
H[176][177]=1;
H[176][353]=1;
H[177][177]=1;
H[177][178]=1;
H[177][270]=3;
H[178][178]=1;
H[178][179]=1;
H[178][319]=1;
H[179][179]=7;
H[179][180]=7;
H[179][376]=1;
H[180][180]=1;
H[180][181]=1;
H[180][345]=1;
H[181][181]=1;
H[181][182]=1;
H[181][308]=1;
H[182][182]=1;
H[182][183]=1;
H[182][338]=1;
H[183][183]=1;
H[183][184]=1;
H[183][327]=1;
H[184][184]=1;
H[184][185]=7;
H[184][273]=7;
H[185][185]=1;
H[185][186]=1;
H[185][381]=1;
H[186][186]=1;
H[186][187]=1;
H[186][299]=2;
H[187][187]=1;
H[187][188]=1;
H[187][280]=1;
H[188][188]=1;
H[188][189]=1;
H[188][357]=1;
H[189][189]=1;
H[189][190]=2;
H[189][292]=1;
H[190][190]=1;
H[190][191]=3;
H[190][311]=1;
H[191][191]=1;
H[191][192]=1;
H[191][341]=2;
H[192][192]=1;
H[192][193]=1;
H[192][349]=1;
H[193][193]=1;
H[193][194]=1;
H[193][370]=6;
H[194][194]=1;
H[194][195]=1;
H[194][321]=3;
H[195][195]=1;
H[195][196]=1;
H[195][282]=1;
H[196][196]=3;
H[196][197]=1;
H[196][335]=1;
H[197][197]=1;
H[197][198]=1;
H[197][306]=2;
H[198][198]=1;
H[198][199]=3;
H[198][295]=3;
H[199][199]=1;
H[199][200]=2;
H[199][373]=1;
H[200][200]=1;
H[200][201]=2;
H[200][287]=1;
H[201][201]=6;
H[201][202]=1;
H[201][364]=1;
H[202][202]=7;
H[202][203]=1;
H[202][340]=6;
H[203][203]=1;
H[203][204]=1;
H[203][318]=1;
H[204][204]=1;
H[204][205]=1;
H[204][382]=1;
H[205][205]=1;
H[205][206]=1;
H[205][304]=1;
H[206][206]=1;
H[206][207]=1;
H[206][360]=7;
H[207][207]=1;
H[207][208]=3;
H[207][375]=3;
H[208][208]=1;
H[208][209]=1;
H[208][313]=1;
H[209][209]=1;
H[209][210]=1;
H[209][298]=3;
H[210][210]=1;
H[210][211]=1;
H[210][368]=1;
H[211][211]=1;
H[211][212]=2;
H[211][286]=1;
H[212][212]=1;
H[212][213]=3;
H[212][323]=1;
H[213][213]=1;
H[213][214]=1;
H[213][383]=7;
H[214][214]=1;
H[214][215]=1;
H[214][309]=1;
H[215][215]=2;
H[215][216]=1;
H[215][331]=1;
H[216][216]=1;
H[216][217]=3;
H[216][348]=1;
H[217][217]=1;
H[217][218]=1;
H[217][296]=1;
H[218][218]=7;
H[218][219]=7;
H[218][377]=1;
H[219][219]=1;
H[219][220]=1;
H[219][284]=1;
H[220][220]=7;
H[220][221]=7;
H[220][358]=1;
H[221][221]=1;
H[221][222]=1;
H[221][328]=1;
H[222][222]=1;
H[222][223]=1;
H[222][372]=1;
H[223][223]=1;
H[223][224]=1;
H[223][276]=1;
H[224][224]=6;
H[224][225]=1;
H[224][301]=1;
H[225][225]=1;
H[225][226]=6;
H[225][316]=7;
H[226][226]=1;
H[226][227]=6;
H[226][332]=1;
H[227][227]=1;
H[227][228]=2;
H[227][380]=1;
H[228][228]=1;
H[228][229]=1;
H[228][291]=1;
H[229][229]=2;
H[229][230]=1;
H[229][362]=1;
H[230][230]=1;
H[230][231]=1;
H[230][283]=1;
H[231][231]=1;
H[231][232]=1;
H[231][274]=1;
H[232][232]=1;
H[232][233]=6;
H[232][346]=1;
H[233][233]=1;
H[233][234]=1;
H[233][354]=2;
H[234][234]=1;
H[234][235]=1;
H[234][333]=1;
H[235][235]=1;
H[235][236]=1;
H[235][369]=1;
H[236][236]=1;
H[236][237]=1;
H[236][263]=1;
H[237][237]=1;
H[237][238]=1;
H[237][361]=1;
H[238][238]=1;
H[238][239]=1;
H[238][271]=1;
H[239][239]=1;
H[239][240]=1;
H[239][310]=2;
H[240][240]=1;
H[240][241]=1;
H[240][379]=1;
H[241][241]=1;
H[241][242]=3;
H[241][366]=3;
H[242][242]=7;
H[242][243]=7;
H[242][281]=1;
H[243][243]=3;
H[243][244]=1;
H[243][260]=3;
H[244][244]=1;
H[244][245]=1;
H[244][317]=1;
H[245][245]=1;
H[245][246]=3;
H[245][347]=1;
H[246][246]=1;
H[246][247]=3;
H[246][267]=1;
H[247][247]=1;
H[247][248]=1;
H[247][290]=1;
H[248][248]=1;
H[248][249]=1;
H[248][303]=3;
H[249][249]=7;
H[249][250]=7;
H[249][365]=1;
H[250][250]=1;
H[250][251]=1;
H[250][329]=1;
H[251][251]=3;
H[251][252]=3;
H[251][258]=1;
H[252][252]=6;
H[252][253]=1;
H[252][352]=7;
H[253][253]=1;
H[253][254]=1;
H[253][312]=1;
H[254][254]=1;
H[254][255]=1;
H[254][275]=1;
H[255][128]=1;
H[255][255]=1;
H[255][324]=1;


/* BELOW IS THE INITIALIZATION FOR THE ROW_COL*/
row_col[0][0]=0;
row_col[1][0]=127;
row_col[0][1]=0;
row_col[1][1]=1;
row_col[0][2]=1;
row_col[1][2]=2;
row_col[0][3]=2;
row_col[1][3]=3;
row_col[0][4]=3;
row_col[1][4]=4;
row_col[0][5]=4;
row_col[1][5]=5;
row_col[0][6]=5;
row_col[1][6]=6;
row_col[0][7]=6;
row_col[1][7]=7;
row_col[0][8]=7;
row_col[1][8]=8;
row_col[0][9]=8;
row_col[1][9]=9;
row_col[0][10]=9;
row_col[1][10]=10;
row_col[0][11]=10;
row_col[1][11]=11;
row_col[0][12]=11;
row_col[1][12]=12;
row_col[0][13]=12;
row_col[1][13]=13;
row_col[0][14]=13;
row_col[1][14]=14;
row_col[0][15]=14;
row_col[1][15]=15;
row_col[0][16]=15;
row_col[1][16]=16;
row_col[0][17]=16;
row_col[1][17]=17;
row_col[0][18]=17;
row_col[1][18]=18;
row_col[0][19]=18;
row_col[1][19]=19;
row_col[0][20]=19;
row_col[1][20]=20;
row_col[0][21]=20;
row_col[1][21]=21;
row_col[0][22]=21;
row_col[1][22]=22;
row_col[0][23]=22;
row_col[1][23]=23;
row_col[0][24]=23;
row_col[1][24]=24;
row_col[0][25]=24;
row_col[1][25]=25;
row_col[0][26]=25;
row_col[1][26]=26;
row_col[0][27]=26;
row_col[1][27]=27;
row_col[0][28]=27;
row_col[1][28]=28;
row_col[0][29]=28;
row_col[1][29]=29;
row_col[0][30]=29;
row_col[1][30]=30;
row_col[0][31]=30;
row_col[1][31]=31;
row_col[0][32]=31;
row_col[1][32]=32;
row_col[0][33]=32;
row_col[1][33]=33;
row_col[0][34]=33;
row_col[1][34]=34;
row_col[0][35]=34;
row_col[1][35]=35;
row_col[0][36]=35;
row_col[1][36]=36;
row_col[0][37]=36;
row_col[1][37]=37;
row_col[0][38]=37;
row_col[1][38]=38;
row_col[0][39]=38;
row_col[1][39]=39;
row_col[0][40]=39;
row_col[1][40]=40;
row_col[0][41]=40;
row_col[1][41]=41;
row_col[0][42]=41;
row_col[1][42]=42;
row_col[0][43]=42;
row_col[1][43]=43;
row_col[0][44]=43;
row_col[1][44]=44;
row_col[0][45]=44;
row_col[1][45]=45;
row_col[0][46]=45;
row_col[1][46]=46;
row_col[0][47]=46;
row_col[1][47]=47;
row_col[0][48]=47;
row_col[1][48]=48;
row_col[0][49]=48;
row_col[1][49]=49;
row_col[0][50]=49;
row_col[1][50]=50;
row_col[0][51]=50;
row_col[1][51]=51;
row_col[0][52]=51;
row_col[1][52]=52;
row_col[0][53]=52;
row_col[1][53]=53;
row_col[0][54]=53;
row_col[1][54]=54;
row_col[0][55]=54;
row_col[1][55]=55;
row_col[0][56]=55;
row_col[1][56]=56;
row_col[0][57]=56;
row_col[1][57]=57;
row_col[0][58]=57;
row_col[1][58]=58;
row_col[0][59]=58;
row_col[1][59]=59;
row_col[0][60]=59;
row_col[1][60]=60;
row_col[0][61]=60;
row_col[1][61]=61;
row_col[0][62]=61;
row_col[1][62]=62;
row_col[0][63]=62;
row_col[1][63]=63;
row_col[0][64]=63;
row_col[1][64]=64;
row_col[0][65]=64;
row_col[1][65]=65;
row_col[0][66]=65;
row_col[1][66]=66;
row_col[0][67]=66;
row_col[1][67]=67;
row_col[0][68]=67;
row_col[1][68]=68;
row_col[0][69]=68;
row_col[1][69]=69;
row_col[0][70]=69;
row_col[1][70]=70;
row_col[0][71]=70;
row_col[1][71]=71;
row_col[0][72]=71;
row_col[1][72]=72;
row_col[0][73]=72;
row_col[1][73]=73;
row_col[0][74]=73;
row_col[1][74]=74;
row_col[0][75]=74;
row_col[1][75]=75;
row_col[0][76]=75;
row_col[1][76]=76;
row_col[0][77]=76;
row_col[1][77]=77;
row_col[0][78]=77;
row_col[1][78]=78;
row_col[0][79]=78;
row_col[1][79]=79;
row_col[0][80]=79;
row_col[1][80]=80;
row_col[0][81]=80;
row_col[1][81]=81;
row_col[0][82]=81;
row_col[1][82]=82;
row_col[0][83]=82;
row_col[1][83]=83;
row_col[0][84]=83;
row_col[1][84]=84;
row_col[0][85]=84;
row_col[1][85]=85;
row_col[0][86]=85;
row_col[1][86]=86;
row_col[0][87]=86;
row_col[1][87]=87;
row_col[0][88]=87;
row_col[1][88]=88;
row_col[0][89]=88;
row_col[1][89]=89;
row_col[0][90]=89;
row_col[1][90]=90;
row_col[0][91]=90;
row_col[1][91]=91;
row_col[0][92]=91;
row_col[1][92]=92;
row_col[0][93]=92;
row_col[1][93]=93;
row_col[0][94]=93;
row_col[1][94]=94;
row_col[0][95]=94;
row_col[1][95]=95;
row_col[0][96]=95;
row_col[1][96]=96;
row_col[0][97]=96;
row_col[1][97]=97;
row_col[0][98]=97;
row_col[1][98]=98;
row_col[0][99]=98;
row_col[1][99]=99;
row_col[0][100]=99;
row_col[1][100]=100;
row_col[0][101]=100;
row_col[1][101]=101;
row_col[0][102]=101;
row_col[1][102]=102;
row_col[0][103]=102;
row_col[1][103]=103;
row_col[0][104]=103;
row_col[1][104]=104;
row_col[0][105]=104;
row_col[1][105]=105;
row_col[0][106]=105;
row_col[1][106]=106;
row_col[0][107]=106;
row_col[1][107]=107;
row_col[0][108]=107;
row_col[1][108]=108;
row_col[0][109]=108;
row_col[1][109]=109;
row_col[0][110]=109;
row_col[1][110]=110;
row_col[0][111]=110;
row_col[1][111]=111;
row_col[0][112]=111;
row_col[1][112]=112;
row_col[0][113]=112;
row_col[1][113]=113;
row_col[0][114]=113;
row_col[1][114]=114;
row_col[0][115]=114;
row_col[1][115]=115;
row_col[0][116]=115;
row_col[1][116]=116;
row_col[0][117]=116;
row_col[1][117]=117;
row_col[0][118]=117;
row_col[1][118]=118;
row_col[0][119]=118;
row_col[1][119]=119;
row_col[0][120]=119;
row_col[1][120]=120;
row_col[0][121]=120;
row_col[1][121]=121;
row_col[0][122]=121;
row_col[1][122]=122;
row_col[0][123]=122;
row_col[1][123]=123;
row_col[0][124]=123;
row_col[1][124]=124;
row_col[0][125]=124;
row_col[1][125]=125;
row_col[0][126]=125;
row_col[1][126]=126;
row_col[0][127]=126;
row_col[1][127]=127;
row_col[0][128]=128;
row_col[1][128]=255;
row_col[0][129]=128;
row_col[1][129]=129;
row_col[0][130]=129;
row_col[1][130]=130;
row_col[0][131]=130;
row_col[1][131]=131;
row_col[0][132]=131;
row_col[1][132]=132;
row_col[0][133]=132;
row_col[1][133]=133;
row_col[0][134]=133;
row_col[1][134]=134;
row_col[0][135]=134;
row_col[1][135]=135;
row_col[0][136]=135;
row_col[1][136]=136;
row_col[0][137]=136;
row_col[1][137]=137;
row_col[0][138]=137;
row_col[1][138]=138;
row_col[0][139]=138;
row_col[1][139]=139;
row_col[0][140]=139;
row_col[1][140]=140;
row_col[0][141]=140;
row_col[1][141]=141;
row_col[0][142]=141;
row_col[1][142]=142;
row_col[0][143]=142;
row_col[1][143]=143;
row_col[0][144]=143;
row_col[1][144]=144;
row_col[0][145]=144;
row_col[1][145]=145;
row_col[0][146]=145;
row_col[1][146]=146;
row_col[0][147]=146;
row_col[1][147]=147;
row_col[0][148]=147;
row_col[1][148]=148;
row_col[0][149]=148;
row_col[1][149]=149;
row_col[0][150]=149;
row_col[1][150]=150;
row_col[0][151]=150;
row_col[1][151]=151;
row_col[0][152]=151;
row_col[1][152]=152;
row_col[0][153]=152;
row_col[1][153]=153;
row_col[0][154]=153;
row_col[1][154]=154;
row_col[0][155]=154;
row_col[1][155]=155;
row_col[0][156]=155;
row_col[1][156]=156;
row_col[0][157]=156;
row_col[1][157]=157;
row_col[0][158]=157;
row_col[1][158]=158;
row_col[0][159]=158;
row_col[1][159]=159;
row_col[0][160]=159;
row_col[1][160]=160;
row_col[0][161]=160;
row_col[1][161]=161;
row_col[0][162]=161;
row_col[1][162]=162;
row_col[0][163]=162;
row_col[1][163]=163;
row_col[0][164]=163;
row_col[1][164]=164;
row_col[0][165]=164;
row_col[1][165]=165;
row_col[0][166]=165;
row_col[1][166]=166;
row_col[0][167]=166;
row_col[1][167]=167;
row_col[0][168]=167;
row_col[1][168]=168;
row_col[0][169]=168;
row_col[1][169]=169;
row_col[0][170]=169;
row_col[1][170]=170;
row_col[0][171]=170;
row_col[1][171]=171;
row_col[0][172]=171;
row_col[1][172]=172;
row_col[0][173]=172;
row_col[1][173]=173;
row_col[0][174]=173;
row_col[1][174]=174;
row_col[0][175]=174;
row_col[1][175]=175;
row_col[0][176]=175;
row_col[1][176]=176;
row_col[0][177]=176;
row_col[1][177]=177;
row_col[0][178]=177;
row_col[1][178]=178;
row_col[0][179]=178;
row_col[1][179]=179;
row_col[0][180]=179;
row_col[1][180]=180;
row_col[0][181]=180;
row_col[1][181]=181;
row_col[0][182]=181;
row_col[1][182]=182;
row_col[0][183]=182;
row_col[1][183]=183;
row_col[0][184]=183;
row_col[1][184]=184;
row_col[0][185]=184;
row_col[1][185]=185;
row_col[0][186]=185;
row_col[1][186]=186;
row_col[0][187]=186;
row_col[1][187]=187;
row_col[0][188]=187;
row_col[1][188]=188;
row_col[0][189]=188;
row_col[1][189]=189;
row_col[0][190]=189;
row_col[1][190]=190;
row_col[0][191]=190;
row_col[1][191]=191;
row_col[0][192]=191;
row_col[1][192]=192;
row_col[0][193]=192;
row_col[1][193]=193;
row_col[0][194]=193;
row_col[1][194]=194;
row_col[0][195]=194;
row_col[1][195]=195;
row_col[0][196]=195;
row_col[1][196]=196;
row_col[0][197]=196;
row_col[1][197]=197;
row_col[0][198]=197;
row_col[1][198]=198;
row_col[0][199]=198;
row_col[1][199]=199;
row_col[0][200]=199;
row_col[1][200]=200;
row_col[0][201]=200;
row_col[1][201]=201;
row_col[0][202]=201;
row_col[1][202]=202;
row_col[0][203]=202;
row_col[1][203]=203;
row_col[0][204]=203;
row_col[1][204]=204;
row_col[0][205]=204;
row_col[1][205]=205;
row_col[0][206]=205;
row_col[1][206]=206;
row_col[0][207]=206;
row_col[1][207]=207;
row_col[0][208]=207;
row_col[1][208]=208;
row_col[0][209]=208;
row_col[1][209]=209;
row_col[0][210]=209;
row_col[1][210]=210;
row_col[0][211]=210;
row_col[1][211]=211;
row_col[0][212]=211;
row_col[1][212]=212;
row_col[0][213]=212;
row_col[1][213]=213;
row_col[0][214]=213;
row_col[1][214]=214;
row_col[0][215]=214;
row_col[1][215]=215;
row_col[0][216]=215;
row_col[1][216]=216;
row_col[0][217]=216;
row_col[1][217]=217;
row_col[0][218]=217;
row_col[1][218]=218;
row_col[0][219]=218;
row_col[1][219]=219;
row_col[0][220]=219;
row_col[1][220]=220;
row_col[0][221]=220;
row_col[1][221]=221;
row_col[0][222]=221;
row_col[1][222]=222;
row_col[0][223]=222;
row_col[1][223]=223;
row_col[0][224]=223;
row_col[1][224]=224;
row_col[0][225]=224;
row_col[1][225]=225;
row_col[0][226]=225;
row_col[1][226]=226;
row_col[0][227]=226;
row_col[1][227]=227;
row_col[0][228]=227;
row_col[1][228]=228;
row_col[0][229]=228;
row_col[1][229]=229;
row_col[0][230]=229;
row_col[1][230]=230;
row_col[0][231]=230;
row_col[1][231]=231;
row_col[0][232]=231;
row_col[1][232]=232;
row_col[0][233]=232;
row_col[1][233]=233;
row_col[0][234]=233;
row_col[1][234]=234;
row_col[0][235]=234;
row_col[1][235]=235;
row_col[0][236]=235;
row_col[1][236]=236;
row_col[0][237]=236;
row_col[1][237]=237;
row_col[0][238]=237;
row_col[1][238]=238;
row_col[0][239]=238;
row_col[1][239]=239;
row_col[0][240]=239;
row_col[1][240]=240;
row_col[0][241]=240;
row_col[1][241]=241;
row_col[0][242]=241;
row_col[1][242]=242;
row_col[0][243]=242;
row_col[1][243]=243;
row_col[0][244]=243;
row_col[1][244]=244;
row_col[0][245]=244;
row_col[1][245]=245;
row_col[0][246]=245;
row_col[1][246]=246;
row_col[0][247]=246;
row_col[1][247]=247;
row_col[0][248]=247;
row_col[1][248]=248;
row_col[0][249]=248;
row_col[1][249]=249;
row_col[0][250]=249;
row_col[1][250]=250;
row_col[0][251]=250;
row_col[1][251]=251;
row_col[0][252]=251;
row_col[1][252]=252;
row_col[0][253]=252;
row_col[1][253]=253;
row_col[0][254]=253;
row_col[1][254]=254;
row_col[0][255]=254;
row_col[1][255]=255;
row_col[0][256]=0;
row_col[1][256]=141;
row_col[0][257]=1;
row_col[1][257]=132;
row_col[0][258]=2;
row_col[1][258]=251;
row_col[0][259]=3;
row_col[1][259]=148;
row_col[0][260]=4;
row_col[1][260]=243;
row_col[0][261]=5;
row_col[1][261]=156;
row_col[0][262]=6;
row_col[1][262]=165;
row_col[0][263]=7;
row_col[1][263]=236;
row_col[0][264]=8;
row_col[1][264]=135;
row_col[0][265]=9;
row_col[1][265]=172;
row_col[0][266]=10;
row_col[1][266]=145;
row_col[0][267]=11;
row_col[1][267]=246;
row_col[0][268]=12;
row_col[1][268]=129;
row_col[0][269]=13;
row_col[1][269]=152;
row_col[0][270]=14;
row_col[1][270]=177;
row_col[0][271]=15;
row_col[1][271]=238;
row_col[0][272]=16;
row_col[1][272]=159;
row_col[0][273]=17;
row_col[1][273]=184;
row_col[0][274]=18;
row_col[1][274]=231;
row_col[0][275]=19;
row_col[1][275]=254;
row_col[0][276]=20;
row_col[1][276]=223;
row_col[0][277]=21;
row_col[1][277]=142;
row_col[0][278]=22;
row_col[1][278]=153;
row_col[0][279]=23;
row_col[1][279]=170;
row_col[0][280]=24;
row_col[1][280]=187;
row_col[0][281]=25;
row_col[1][281]=242;
row_col[0][282]=26;
row_col[1][282]=195;
row_col[0][283]=27;
row_col[1][283]=230;
row_col[0][284]=28;
row_col[1][284]=219;
row_col[0][285]=29;
row_col[1][285]=174;
row_col[0][286]=30;
row_col[1][286]=211;
row_col[0][287]=31;
row_col[1][287]=200;
row_col[0][288]=32;
row_col[1][288]=167;
row_col[0][289]=33;
row_col[1][289]=138;
row_col[0][290]=34;
row_col[1][290]=247;
row_col[0][291]=35;
row_col[1][291]=228;
row_col[0][292]=36;
row_col[1][292]=189;
row_col[0][293]=37;
row_col[1][293]=150;
row_col[0][294]=38;
row_col[1][294]=163;
row_col[0][295]=39;
row_col[1][295]=198;
row_col[0][296]=40;
row_col[1][296]=217;
row_col[0][297]=41;
row_col[1][297]=134;
row_col[0][298]=42;
row_col[1][298]=209;
row_col[0][299]=43;
row_col[1][299]=186;
row_col[0][300]=44;
row_col[1][300]=147;
row_col[0][301]=45;
row_col[1][301]=224;
row_col[0][302]=46;
row_col[1][302]=175;
row_col[0][303]=47;
row_col[1][303]=248;
row_col[0][304]=48;
row_col[1][304]=205;
row_col[0][305]=49;
row_col[1][305]=158;
row_col[0][306]=50;
row_col[1][306]=197;
row_col[0][307]=51;
row_col[1][307]=144;
row_col[0][308]=52;
row_col[1][308]=181;
row_col[0][309]=53;
row_col[1][309]=214;
row_col[0][310]=54;
row_col[1][310]=239;
row_col[0][311]=55;
row_col[1][311]=190;
row_col[0][312]=56;
row_col[1][312]=253;
row_col[0][313]=57;
row_col[1][313]=208;
row_col[0][314]=58;
row_col[1][314]=139;
row_col[0][315]=59;
row_col[1][315]=162;
row_col[0][316]=60;
row_col[1][316]=225;
row_col[0][317]=61;
row_col[1][317]=244;
row_col[0][318]=62;
row_col[1][318]=203;
row_col[0][319]=63;
row_col[1][319]=178;
row_col[0][320]=64;
row_col[1][320]=133;
row_col[0][321]=65;
row_col[1][321]=194;
row_col[0][322]=66;
row_col[1][322]=155;
row_col[0][323]=67;
row_col[1][323]=212;
row_col[0][324]=68;
row_col[1][324]=255;
row_col[0][325]=69;
row_col[1][325]=149;
row_col[0][326]=70;
row_col[1][326]=136;
row_col[0][327]=71;
row_col[1][327]=183;
row_col[0][328]=72;
row_col[1][328]=221;
row_col[0][329]=73;
row_col[1][329]=250;
row_col[0][330]=74;
row_col[1][330]=168;
row_col[0][331]=75;
row_col[1][331]=215;
row_col[0][332]=76;
row_col[1][332]=226;
row_col[0][333]=77;
row_col[1][333]=234;
row_col[0][334]=78;
row_col[1][334]=128;
row_col[0][335]=79;
row_col[1][335]=196;
row_col[0][336]=80;
row_col[1][336]=140;
row_col[0][337]=81;
row_col[1][337]=173;
row_col[0][338]=82;
row_col[1][338]=182;
row_col[0][339]=83;
row_col[1][339]=154;
row_col[0][340]=84;
row_col[1][340]=202;
row_col[0][341]=85;
row_col[1][341]=191;
row_col[0][342]=86;
row_col[1][342]=131;
row_col[0][343]=87;
row_col[1][343]=169;
row_col[0][344]=88;
row_col[1][344]=161;
row_col[0][345]=89;
row_col[1][345]=180;
row_col[0][346]=90;
row_col[1][346]=232;
row_col[0][347]=91;
row_col[1][347]=245;
row_col[0][348]=92;
row_col[1][348]=216;
row_col[0][349]=93;
row_col[1][349]=192;
row_col[0][350]=94;
row_col[1][350]=143;
row_col[0][351]=95;
row_col[1][351]=164;
row_col[0][352]=96;
row_col[1][352]=252;
row_col[0][353]=97;
row_col[1][353]=176;
row_col[0][354]=98;
row_col[1][354]=233;
row_col[0][355]=99;
row_col[1][355]=137;
row_col[0][356]=100;
row_col[1][356]=157;
row_col[0][357]=101;
row_col[1][357]=188;
row_col[0][358]=102;
row_col[1][358]=220;
row_col[0][359]=103;
row_col[1][359]=130;
row_col[0][360]=104;
row_col[1][360]=206;
row_col[0][361]=105;
row_col[1][361]=237;
row_col[0][362]=106;
row_col[1][362]=229;
row_col[0][363]=107;
row_col[1][363]=146;
row_col[0][364]=108;
row_col[1][364]=201;
row_col[0][365]=109;
row_col[1][365]=249;
row_col[0][366]=110;
row_col[1][366]=241;
row_col[0][367]=111;
row_col[1][367]=151;
row_col[0][368]=112;
row_col[1][368]=210;
row_col[0][369]=113;
row_col[1][369]=235;
row_col[0][370]=114;
row_col[1][370]=193;
row_col[0][371]=115;
row_col[1][371]=160;
row_col[0][372]=116;
row_col[1][372]=222;
row_col[0][373]=117;
row_col[1][373]=199;
row_col[0][374]=118;
row_col[1][374]=171;
row_col[0][375]=119;
row_col[1][375]=207;
row_col[0][376]=120;
row_col[1][376]=179;
row_col[0][377]=121;
row_col[1][377]=218;
row_col[0][378]=122;
row_col[1][378]=166;
row_col[0][379]=123;
row_col[1][379]=240;
row_col[0][380]=124;
row_col[1][380]=227;
row_col[0][381]=125;
row_col[1][381]=185;
row_col[0][382]=126;
row_col[1][382]=204;
row_col[0][383]=127;
row_col[1][383]=213;

/*BELOW IS THE INITIALIZATION FOR COL_ROW*/
col_row[0][0]=0;
col_row[0][1]=1;
col_row[0][2]=256;
col_row[1][0]=1;
col_row[1][1]=2;
col_row[1][2]=257;
col_row[2][0]=2;
col_row[2][1]=3;
col_row[2][2]=258;
col_row[3][0]=3;
col_row[3][1]=4;
col_row[3][2]=259;
col_row[4][0]=4;
col_row[4][1]=5;
col_row[4][2]=260;
col_row[5][0]=5;
col_row[5][1]=6;
col_row[5][2]=261;
col_row[6][0]=6;
col_row[6][1]=7;
col_row[6][2]=262;
col_row[7][0]=7;
col_row[7][1]=8;
col_row[7][2]=263;
col_row[8][0]=8;
col_row[8][1]=9;
col_row[8][2]=264;
col_row[9][0]=9;
col_row[9][1]=10;
col_row[9][2]=265;
col_row[10][0]=10;
col_row[10][1]=11;
col_row[10][2]=266;
col_row[11][0]=11;
col_row[11][1]=12;
col_row[11][2]=267;
col_row[12][0]=12;
col_row[12][1]=13;
col_row[12][2]=268;
col_row[13][0]=13;
col_row[13][1]=14;
col_row[13][2]=269;
col_row[14][0]=14;
col_row[14][1]=15;
col_row[14][2]=270;
col_row[15][0]=15;
col_row[15][1]=16;
col_row[15][2]=271;
col_row[16][0]=16;
col_row[16][1]=17;
col_row[16][2]=272;
col_row[17][0]=17;
col_row[17][1]=18;
col_row[17][2]=273;
col_row[18][0]=18;
col_row[18][1]=19;
col_row[18][2]=274;
col_row[19][0]=19;
col_row[19][1]=20;
col_row[19][2]=275;
col_row[20][0]=20;
col_row[20][1]=21;
col_row[20][2]=276;
col_row[21][0]=21;
col_row[21][1]=22;
col_row[21][2]=277;
col_row[22][0]=22;
col_row[22][1]=23;
col_row[22][2]=278;
col_row[23][0]=23;
col_row[23][1]=24;
col_row[23][2]=279;
col_row[24][0]=24;
col_row[24][1]=25;
col_row[24][2]=280;
col_row[25][0]=25;
col_row[25][1]=26;
col_row[25][2]=281;
col_row[26][0]=26;
col_row[26][1]=27;
col_row[26][2]=282;
col_row[27][0]=27;
col_row[27][1]=28;
col_row[27][2]=283;
col_row[28][0]=28;
col_row[28][1]=29;
col_row[28][2]=284;
col_row[29][0]=29;
col_row[29][1]=30;
col_row[29][2]=285;
col_row[30][0]=30;
col_row[30][1]=31;
col_row[30][2]=286;
col_row[31][0]=31;
col_row[31][1]=32;
col_row[31][2]=287;
col_row[32][0]=32;
col_row[32][1]=33;
col_row[32][2]=288;
col_row[33][0]=33;
col_row[33][1]=34;
col_row[33][2]=289;
col_row[34][0]=34;
col_row[34][1]=35;
col_row[34][2]=290;
col_row[35][0]=35;
col_row[35][1]=36;
col_row[35][2]=291;
col_row[36][0]=36;
col_row[36][1]=37;
col_row[36][2]=292;
col_row[37][0]=37;
col_row[37][1]=38;
col_row[37][2]=293;
col_row[38][0]=38;
col_row[38][1]=39;
col_row[38][2]=294;
col_row[39][0]=39;
col_row[39][1]=40;
col_row[39][2]=295;
col_row[40][0]=40;
col_row[40][1]=41;
col_row[40][2]=296;
col_row[41][0]=41;
col_row[41][1]=42;
col_row[41][2]=297;
col_row[42][0]=42;
col_row[42][1]=43;
col_row[42][2]=298;
col_row[43][0]=43;
col_row[43][1]=44;
col_row[43][2]=299;
col_row[44][0]=44;
col_row[44][1]=45;
col_row[44][2]=300;
col_row[45][0]=45;
col_row[45][1]=46;
col_row[45][2]=301;
col_row[46][0]=46;
col_row[46][1]=47;
col_row[46][2]=302;
col_row[47][0]=47;
col_row[47][1]=48;
col_row[47][2]=303;
col_row[48][0]=48;
col_row[48][1]=49;
col_row[48][2]=304;
col_row[49][0]=49;
col_row[49][1]=50;
col_row[49][2]=305;
col_row[50][0]=50;
col_row[50][1]=51;
col_row[50][2]=306;
col_row[51][0]=51;
col_row[51][1]=52;
col_row[51][2]=307;
col_row[52][0]=52;
col_row[52][1]=53;
col_row[52][2]=308;
col_row[53][0]=53;
col_row[53][1]=54;
col_row[53][2]=309;
col_row[54][0]=54;
col_row[54][1]=55;
col_row[54][2]=310;
col_row[55][0]=55;
col_row[55][1]=56;
col_row[55][2]=311;
col_row[56][0]=56;
col_row[56][1]=57;
col_row[56][2]=312;
col_row[57][0]=57;
col_row[57][1]=58;
col_row[57][2]=313;
col_row[58][0]=58;
col_row[58][1]=59;
col_row[58][2]=314;
col_row[59][0]=59;
col_row[59][1]=60;
col_row[59][2]=315;
col_row[60][0]=60;
col_row[60][1]=61;
col_row[60][2]=316;
col_row[61][0]=61;
col_row[61][1]=62;
col_row[61][2]=317;
col_row[62][0]=62;
col_row[62][1]=63;
col_row[62][2]=318;
col_row[63][0]=63;
col_row[63][1]=64;
col_row[63][2]=319;
col_row[64][0]=64;
col_row[64][1]=65;
col_row[64][2]=320;
col_row[65][0]=65;
col_row[65][1]=66;
col_row[65][2]=321;
col_row[66][0]=66;
col_row[66][1]=67;
col_row[66][2]=322;
col_row[67][0]=67;
col_row[67][1]=68;
col_row[67][2]=323;
col_row[68][0]=68;
col_row[68][1]=69;
col_row[68][2]=324;
col_row[69][0]=69;
col_row[69][1]=70;
col_row[69][2]=325;
col_row[70][0]=70;
col_row[70][1]=71;
col_row[70][2]=326;
col_row[71][0]=71;
col_row[71][1]=72;
col_row[71][2]=327;
col_row[72][0]=72;
col_row[72][1]=73;
col_row[72][2]=328;
col_row[73][0]=73;
col_row[73][1]=74;
col_row[73][2]=329;
col_row[74][0]=74;
col_row[74][1]=75;
col_row[74][2]=330;
col_row[75][0]=75;
col_row[75][1]=76;
col_row[75][2]=331;
col_row[76][0]=76;
col_row[76][1]=77;
col_row[76][2]=332;
col_row[77][0]=77;
col_row[77][1]=78;
col_row[77][2]=333;
col_row[78][0]=78;
col_row[78][1]=79;
col_row[78][2]=334;
col_row[79][0]=79;
col_row[79][1]=80;
col_row[79][2]=335;
col_row[80][0]=80;
col_row[80][1]=81;
col_row[80][2]=336;
col_row[81][0]=81;
col_row[81][1]=82;
col_row[81][2]=337;
col_row[82][0]=82;
col_row[82][1]=83;
col_row[82][2]=338;
col_row[83][0]=83;
col_row[83][1]=84;
col_row[83][2]=339;
col_row[84][0]=84;
col_row[84][1]=85;
col_row[84][2]=340;
col_row[85][0]=85;
col_row[85][1]=86;
col_row[85][2]=341;
col_row[86][0]=86;
col_row[86][1]=87;
col_row[86][2]=342;
col_row[87][0]=87;
col_row[87][1]=88;
col_row[87][2]=343;
col_row[88][0]=88;
col_row[88][1]=89;
col_row[88][2]=344;
col_row[89][0]=89;
col_row[89][1]=90;
col_row[89][2]=345;
col_row[90][0]=90;
col_row[90][1]=91;
col_row[90][2]=346;
col_row[91][0]=91;
col_row[91][1]=92;
col_row[91][2]=347;
col_row[92][0]=92;
col_row[92][1]=93;
col_row[92][2]=348;
col_row[93][0]=93;
col_row[93][1]=94;
col_row[93][2]=349;
col_row[94][0]=94;
col_row[94][1]=95;
col_row[94][2]=350;
col_row[95][0]=95;
col_row[95][1]=96;
col_row[95][2]=351;
col_row[96][0]=96;
col_row[96][1]=97;
col_row[96][2]=352;
col_row[97][0]=97;
col_row[97][1]=98;
col_row[97][2]=353;
col_row[98][0]=98;
col_row[98][1]=99;
col_row[98][2]=354;
col_row[99][0]=99;
col_row[99][1]=100;
col_row[99][2]=355;
col_row[100][0]=100;
col_row[100][1]=101;
col_row[100][2]=356;
col_row[101][0]=101;
col_row[101][1]=102;
col_row[101][2]=357;
col_row[102][0]=102;
col_row[102][1]=103;
col_row[102][2]=358;
col_row[103][0]=103;
col_row[103][1]=104;
col_row[103][2]=359;
col_row[104][0]=104;
col_row[104][1]=105;
col_row[104][2]=360;
col_row[105][0]=105;
col_row[105][1]=106;
col_row[105][2]=361;
col_row[106][0]=106;
col_row[106][1]=107;
col_row[106][2]=362;
col_row[107][0]=107;
col_row[107][1]=108;
col_row[107][2]=363;
col_row[108][0]=108;
col_row[108][1]=109;
col_row[108][2]=364;
col_row[109][0]=109;
col_row[109][1]=110;
col_row[109][2]=365;
col_row[110][0]=110;
col_row[110][1]=111;
col_row[110][2]=366;
col_row[111][0]=111;
col_row[111][1]=112;
col_row[111][2]=367;
col_row[112][0]=112;
col_row[112][1]=113;
col_row[112][2]=368;
col_row[113][0]=113;
col_row[113][1]=114;
col_row[113][2]=369;
col_row[114][0]=114;
col_row[114][1]=115;
col_row[114][2]=370;
col_row[115][0]=115;
col_row[115][1]=116;
col_row[115][2]=371;
col_row[116][0]=116;
col_row[116][1]=117;
col_row[116][2]=372;
col_row[117][0]=117;
col_row[117][1]=118;
col_row[117][2]=373;
col_row[118][0]=118;
col_row[118][1]=119;
col_row[118][2]=374;
col_row[119][0]=119;
col_row[119][1]=120;
col_row[119][2]=375;
col_row[120][0]=120;
col_row[120][1]=121;
col_row[120][2]=376;
col_row[121][0]=121;
col_row[121][1]=122;
col_row[121][2]=377;
col_row[122][0]=122;
col_row[122][1]=123;
col_row[122][2]=378;
col_row[123][0]=123;
col_row[123][1]=124;
col_row[123][2]=379;
col_row[124][0]=124;
col_row[124][1]=125;
col_row[124][2]=380;
col_row[125][0]=125;
col_row[125][1]=126;
col_row[125][2]=381;
col_row[126][0]=126;
col_row[126][1]=127;
col_row[126][2]=382;
col_row[127][0]=0;
col_row[127][1]=127;
col_row[127][2]=383;
col_row[128][0]=128;
col_row[128][1]=129;
col_row[128][2]=334;
col_row[129][0]=129;
col_row[129][1]=130;
col_row[129][2]=268;
col_row[130][0]=130;
col_row[130][1]=131;
col_row[130][2]=359;
col_row[131][0]=131;
col_row[131][1]=132;
col_row[131][2]=342;
col_row[132][0]=132;
col_row[132][1]=133;
col_row[132][2]=257;
col_row[133][0]=133;
col_row[133][1]=134;
col_row[133][2]=320;
col_row[134][0]=134;
col_row[134][1]=135;
col_row[134][2]=297;
col_row[135][0]=135;
col_row[135][1]=136;
col_row[135][2]=264;
col_row[136][0]=136;
col_row[136][1]=137;
col_row[136][2]=326;
col_row[137][0]=137;
col_row[137][1]=138;
col_row[137][2]=355;
col_row[138][0]=138;
col_row[138][1]=139;
col_row[138][2]=289;
col_row[139][0]=139;
col_row[139][1]=140;
col_row[139][2]=314;
col_row[140][0]=140;
col_row[140][1]=141;
col_row[140][2]=336;
col_row[141][0]=141;
col_row[141][1]=142;
col_row[141][2]=256;
col_row[142][0]=142;
col_row[142][1]=143;
col_row[142][2]=277;
col_row[143][0]=143;
col_row[143][1]=144;
col_row[143][2]=350;
col_row[144][0]=144;
col_row[144][1]=145;
col_row[144][2]=307;
col_row[145][0]=145;
col_row[145][1]=146;
col_row[145][2]=266;
col_row[146][0]=146;
col_row[146][1]=147;
col_row[146][2]=363;
col_row[147][0]=147;
col_row[147][1]=148;
col_row[147][2]=300;
col_row[148][0]=148;
col_row[148][1]=149;
col_row[148][2]=259;
col_row[149][0]=149;
col_row[149][1]=150;
col_row[149][2]=325;
col_row[150][0]=150;
col_row[150][1]=151;
col_row[150][2]=293;
col_row[151][0]=151;
col_row[151][1]=152;
col_row[151][2]=367;
col_row[152][0]=152;
col_row[152][1]=153;
col_row[152][2]=269;
col_row[153][0]=153;
col_row[153][1]=154;
col_row[153][2]=278;
col_row[154][0]=154;
col_row[154][1]=155;
col_row[154][2]=339;
col_row[155][0]=155;
col_row[155][1]=156;
col_row[155][2]=322;
col_row[156][0]=156;
col_row[156][1]=157;
col_row[156][2]=261;
col_row[157][0]=157;
col_row[157][1]=158;
col_row[157][2]=356;
col_row[158][0]=158;
col_row[158][1]=159;
col_row[158][2]=305;
col_row[159][0]=159;
col_row[159][1]=160;
col_row[159][2]=272;
col_row[160][0]=160;
col_row[160][1]=161;
col_row[160][2]=371;
col_row[161][0]=161;
col_row[161][1]=162;
col_row[161][2]=344;
col_row[162][0]=162;
col_row[162][1]=163;
col_row[162][2]=315;
col_row[163][0]=163;
col_row[163][1]=164;
col_row[163][2]=294;
col_row[164][0]=164;
col_row[164][1]=165;
col_row[164][2]=351;
col_row[165][0]=165;
col_row[165][1]=166;
col_row[165][2]=262;
col_row[166][0]=166;
col_row[166][1]=167;
col_row[166][2]=378;
col_row[167][0]=167;
col_row[167][1]=168;
col_row[167][2]=288;
col_row[168][0]=168;
col_row[168][1]=169;
col_row[168][2]=330;
col_row[169][0]=169;
col_row[169][1]=170;
col_row[169][2]=343;
col_row[170][0]=170;
col_row[170][1]=171;
col_row[170][2]=279;
col_row[171][0]=171;
col_row[171][1]=172;
col_row[171][2]=374;
col_row[172][0]=172;
col_row[172][1]=173;
col_row[172][2]=265;
col_row[173][0]=173;
col_row[173][1]=174;
col_row[173][2]=337;
col_row[174][0]=174;
col_row[174][1]=175;
col_row[174][2]=285;
col_row[175][0]=175;
col_row[175][1]=176;
col_row[175][2]=302;
col_row[176][0]=176;
col_row[176][1]=177;
col_row[176][2]=353;
col_row[177][0]=177;
col_row[177][1]=178;
col_row[177][2]=270;
col_row[178][0]=178;
col_row[178][1]=179;
col_row[178][2]=319;
col_row[179][0]=179;
col_row[179][1]=180;
col_row[179][2]=376;
col_row[180][0]=180;
col_row[180][1]=181;
col_row[180][2]=345;
col_row[181][0]=181;
col_row[181][1]=182;
col_row[181][2]=308;
col_row[182][0]=182;
col_row[182][1]=183;
col_row[182][2]=338;
col_row[183][0]=183;
col_row[183][1]=184;
col_row[183][2]=327;
col_row[184][0]=184;
col_row[184][1]=185;
col_row[184][2]=273;
col_row[185][0]=185;
col_row[185][1]=186;
col_row[185][2]=381;
col_row[186][0]=186;
col_row[186][1]=187;
col_row[186][2]=299;
col_row[187][0]=187;
col_row[187][1]=188;
col_row[187][2]=280;
col_row[188][0]=188;
col_row[188][1]=189;
col_row[188][2]=357;
col_row[189][0]=189;
col_row[189][1]=190;
col_row[189][2]=292;
col_row[190][0]=190;
col_row[190][1]=191;
col_row[190][2]=311;
col_row[191][0]=191;
col_row[191][1]=192;
col_row[191][2]=341;
col_row[192][0]=192;
col_row[192][1]=193;
col_row[192][2]=349;
col_row[193][0]=193;
col_row[193][1]=194;
col_row[193][2]=370;
col_row[194][0]=194;
col_row[194][1]=195;
col_row[194][2]=321;
col_row[195][0]=195;
col_row[195][1]=196;
col_row[195][2]=282;
col_row[196][0]=196;
col_row[196][1]=197;
col_row[196][2]=335;
col_row[197][0]=197;
col_row[197][1]=198;
col_row[197][2]=306;
col_row[198][0]=198;
col_row[198][1]=199;
col_row[198][2]=295;
col_row[199][0]=199;
col_row[199][1]=200;
col_row[199][2]=373;
col_row[200][0]=200;
col_row[200][1]=201;
col_row[200][2]=287;
col_row[201][0]=201;
col_row[201][1]=202;
col_row[201][2]=364;
col_row[202][0]=202;
col_row[202][1]=203;
col_row[202][2]=340;
col_row[203][0]=203;
col_row[203][1]=204;
col_row[203][2]=318;
col_row[204][0]=204;
col_row[204][1]=205;
col_row[204][2]=382;
col_row[205][0]=205;
col_row[205][1]=206;
col_row[205][2]=304;
col_row[206][0]=206;
col_row[206][1]=207;
col_row[206][2]=360;
col_row[207][0]=207;
col_row[207][1]=208;
col_row[207][2]=375;
col_row[208][0]=208;
col_row[208][1]=209;
col_row[208][2]=313;
col_row[209][0]=209;
col_row[209][1]=210;
col_row[209][2]=298;
col_row[210][0]=210;
col_row[210][1]=211;
col_row[210][2]=368;
col_row[211][0]=211;
col_row[211][1]=212;
col_row[211][2]=286;
col_row[212][0]=212;
col_row[212][1]=213;
col_row[212][2]=323;
col_row[213][0]=213;
col_row[213][1]=214;
col_row[213][2]=383;
col_row[214][0]=214;
col_row[214][1]=215;
col_row[214][2]=309;
col_row[215][0]=215;
col_row[215][1]=216;
col_row[215][2]=331;
col_row[216][0]=216;
col_row[216][1]=217;
col_row[216][2]=348;
col_row[217][0]=217;
col_row[217][1]=218;
col_row[217][2]=296;
col_row[218][0]=218;
col_row[218][1]=219;
col_row[218][2]=377;
col_row[219][0]=219;
col_row[219][1]=220;
col_row[219][2]=284;
col_row[220][0]=220;
col_row[220][1]=221;
col_row[220][2]=358;
col_row[221][0]=221;
col_row[221][1]=222;
col_row[221][2]=328;
col_row[222][0]=222;
col_row[222][1]=223;
col_row[222][2]=372;
col_row[223][0]=223;
col_row[223][1]=224;
col_row[223][2]=276;
col_row[224][0]=224;
col_row[224][1]=225;
col_row[224][2]=301;
col_row[225][0]=225;
col_row[225][1]=226;
col_row[225][2]=316;
col_row[226][0]=226;
col_row[226][1]=227;
col_row[226][2]=332;
col_row[227][0]=227;
col_row[227][1]=228;
col_row[227][2]=380;
col_row[228][0]=228;
col_row[228][1]=229;
col_row[228][2]=291;
col_row[229][0]=229;
col_row[229][1]=230;
col_row[229][2]=362;
col_row[230][0]=230;
col_row[230][1]=231;
col_row[230][2]=283;
col_row[231][0]=231;
col_row[231][1]=232;
col_row[231][2]=274;
col_row[232][0]=232;
col_row[232][1]=233;
col_row[232][2]=346;
col_row[233][0]=233;
col_row[233][1]=234;
col_row[233][2]=354;
col_row[234][0]=234;
col_row[234][1]=235;
col_row[234][2]=333;
col_row[235][0]=235;
col_row[235][1]=236;
col_row[235][2]=369;
col_row[236][0]=236;
col_row[236][1]=237;
col_row[236][2]=263;
col_row[237][0]=237;
col_row[237][1]=238;
col_row[237][2]=361;
col_row[238][0]=238;
col_row[238][1]=239;
col_row[238][2]=271;
col_row[239][0]=239;
col_row[239][1]=240;
col_row[239][2]=310;
col_row[240][0]=240;
col_row[240][1]=241;
col_row[240][2]=379;
col_row[241][0]=241;
col_row[241][1]=242;
col_row[241][2]=366;
col_row[242][0]=242;
col_row[242][1]=243;
col_row[242][2]=281;
col_row[243][0]=243;
col_row[243][1]=244;
col_row[243][2]=260;
col_row[244][0]=244;
col_row[244][1]=245;
col_row[244][2]=317;
col_row[245][0]=245;
col_row[245][1]=246;
col_row[245][2]=347;
col_row[246][0]=246;
col_row[246][1]=247;
col_row[246][2]=267;
col_row[247][0]=247;
col_row[247][1]=248;
col_row[247][2]=290;
col_row[248][0]=248;
col_row[248][1]=249;
col_row[248][2]=303;
col_row[249][0]=249;
col_row[249][1]=250;
col_row[249][2]=365;
col_row[250][0]=250;
col_row[250][1]=251;
col_row[250][2]=329;
col_row[251][0]=251;
col_row[251][1]=252;
col_row[251][2]=258;
col_row[252][0]=252;
col_row[252][1]=253;
col_row[252][2]=352;
col_row[253][0]=253;
col_row[253][1]=254;
col_row[253][2]=312;
col_row[254][0]=254;
col_row[254][1]=255;
col_row[254][2]=275;
col_row[255][0]=128;
col_row[255][1]=255;
col_row[255][2]=324;

/* BELOW IS THE INITIALIZATION FOR MAGICV*/
index_VN[0][0]=0;
index_VN[127][0]=1;
index_VN[0][1]=0;
index_VN[1][1]=1;
index_VN[1][2]=0;
index_VN[2][2]=1;
index_VN[2][3]=0;
index_VN[3][3]=1;
index_VN[3][4]=0;
index_VN[4][4]=1;
index_VN[4][5]=0;
index_VN[5][5]=1;
index_VN[5][6]=0;
index_VN[6][6]=1;
index_VN[6][7]=0;
index_VN[7][7]=1;
index_VN[7][8]=0;
index_VN[8][8]=1;
index_VN[8][9]=0;
index_VN[9][9]=1;
index_VN[9][10]=0;
index_VN[10][10]=1;
index_VN[10][11]=0;
index_VN[11][11]=1;
index_VN[11][12]=0;
index_VN[12][12]=1;
index_VN[12][13]=0;
index_VN[13][13]=1;
index_VN[13][14]=0;
index_VN[14][14]=1;
index_VN[14][15]=0;
index_VN[15][15]=1;
index_VN[15][16]=0;
index_VN[16][16]=1;
index_VN[16][17]=0;
index_VN[17][17]=1;
index_VN[17][18]=0;
index_VN[18][18]=1;
index_VN[18][19]=0;
index_VN[19][19]=1;
index_VN[19][20]=0;
index_VN[20][20]=1;
index_VN[20][21]=0;
index_VN[21][21]=1;
index_VN[21][22]=0;
index_VN[22][22]=1;
index_VN[22][23]=0;
index_VN[23][23]=1;
index_VN[23][24]=0;
index_VN[24][24]=1;
index_VN[24][25]=0;
index_VN[25][25]=1;
index_VN[25][26]=0;
index_VN[26][26]=1;
index_VN[26][27]=0;
index_VN[27][27]=1;
index_VN[27][28]=0;
index_VN[28][28]=1;
index_VN[28][29]=0;
index_VN[29][29]=1;
index_VN[29][30]=0;
index_VN[30][30]=1;
index_VN[30][31]=0;
index_VN[31][31]=1;
index_VN[31][32]=0;
index_VN[32][32]=1;
index_VN[32][33]=0;
index_VN[33][33]=1;
index_VN[33][34]=0;
index_VN[34][34]=1;
index_VN[34][35]=0;
index_VN[35][35]=1;
index_VN[35][36]=0;
index_VN[36][36]=1;
index_VN[36][37]=0;
index_VN[37][37]=1;
index_VN[37][38]=0;
index_VN[38][38]=1;
index_VN[38][39]=0;
index_VN[39][39]=1;
index_VN[39][40]=0;
index_VN[40][40]=1;
index_VN[40][41]=0;
index_VN[41][41]=1;
index_VN[41][42]=0;
index_VN[42][42]=1;
index_VN[42][43]=0;
index_VN[43][43]=1;
index_VN[43][44]=0;
index_VN[44][44]=1;
index_VN[44][45]=0;
index_VN[45][45]=1;
index_VN[45][46]=0;
index_VN[46][46]=1;
index_VN[46][47]=0;
index_VN[47][47]=1;
index_VN[47][48]=0;
index_VN[48][48]=1;
index_VN[48][49]=0;
index_VN[49][49]=1;
index_VN[49][50]=0;
index_VN[50][50]=1;
index_VN[50][51]=0;
index_VN[51][51]=1;
index_VN[51][52]=0;
index_VN[52][52]=1;
index_VN[52][53]=0;
index_VN[53][53]=1;
index_VN[53][54]=0;
index_VN[54][54]=1;
index_VN[54][55]=0;
index_VN[55][55]=1;
index_VN[55][56]=0;
index_VN[56][56]=1;
index_VN[56][57]=0;
index_VN[57][57]=1;
index_VN[57][58]=0;
index_VN[58][58]=1;
index_VN[58][59]=0;
index_VN[59][59]=1;
index_VN[59][60]=0;
index_VN[60][60]=1;
index_VN[60][61]=0;
index_VN[61][61]=1;
index_VN[61][62]=0;
index_VN[62][62]=1;
index_VN[62][63]=0;
index_VN[63][63]=1;
index_VN[63][64]=0;
index_VN[64][64]=1;
index_VN[64][65]=0;
index_VN[65][65]=1;
index_VN[65][66]=0;
index_VN[66][66]=1;
index_VN[66][67]=0;
index_VN[67][67]=1;
index_VN[67][68]=0;
index_VN[68][68]=1;
index_VN[68][69]=0;
index_VN[69][69]=1;
index_VN[69][70]=0;
index_VN[70][70]=1;
index_VN[70][71]=0;
index_VN[71][71]=1;
index_VN[71][72]=0;
index_VN[72][72]=1;
index_VN[72][73]=0;
index_VN[73][73]=1;
index_VN[73][74]=0;
index_VN[74][74]=1;
index_VN[74][75]=0;
index_VN[75][75]=1;
index_VN[75][76]=0;
index_VN[76][76]=1;
index_VN[76][77]=0;
index_VN[77][77]=1;
index_VN[77][78]=0;
index_VN[78][78]=1;
index_VN[78][79]=0;
index_VN[79][79]=1;
index_VN[79][80]=0;
index_VN[80][80]=1;
index_VN[80][81]=0;
index_VN[81][81]=1;
index_VN[81][82]=0;
index_VN[82][82]=1;
index_VN[82][83]=0;
index_VN[83][83]=1;
index_VN[83][84]=0;
index_VN[84][84]=1;
index_VN[84][85]=0;
index_VN[85][85]=1;
index_VN[85][86]=0;
index_VN[86][86]=1;
index_VN[86][87]=0;
index_VN[87][87]=1;
index_VN[87][88]=0;
index_VN[88][88]=1;
index_VN[88][89]=0;
index_VN[89][89]=1;
index_VN[89][90]=0;
index_VN[90][90]=1;
index_VN[90][91]=0;
index_VN[91][91]=1;
index_VN[91][92]=0;
index_VN[92][92]=1;
index_VN[92][93]=0;
index_VN[93][93]=1;
index_VN[93][94]=0;
index_VN[94][94]=1;
index_VN[94][95]=0;
index_VN[95][95]=1;
index_VN[95][96]=0;
index_VN[96][96]=1;
index_VN[96][97]=0;
index_VN[97][97]=1;
index_VN[97][98]=0;
index_VN[98][98]=1;
index_VN[98][99]=0;
index_VN[99][99]=1;
index_VN[99][100]=0;
index_VN[100][100]=1;
index_VN[100][101]=0;
index_VN[101][101]=1;
index_VN[101][102]=0;
index_VN[102][102]=1;
index_VN[102][103]=0;
index_VN[103][103]=1;
index_VN[103][104]=0;
index_VN[104][104]=1;
index_VN[104][105]=0;
index_VN[105][105]=1;
index_VN[105][106]=0;
index_VN[106][106]=1;
index_VN[106][107]=0;
index_VN[107][107]=1;
index_VN[107][108]=0;
index_VN[108][108]=1;
index_VN[108][109]=0;
index_VN[109][109]=1;
index_VN[109][110]=0;
index_VN[110][110]=1;
index_VN[110][111]=0;
index_VN[111][111]=1;
index_VN[111][112]=0;
index_VN[112][112]=1;
index_VN[112][113]=0;
index_VN[113][113]=1;
index_VN[113][114]=0;
index_VN[114][114]=1;
index_VN[114][115]=0;
index_VN[115][115]=1;
index_VN[115][116]=0;
index_VN[116][116]=1;
index_VN[116][117]=0;
index_VN[117][117]=1;
index_VN[117][118]=0;
index_VN[118][118]=1;
index_VN[118][119]=0;
index_VN[119][119]=1;
index_VN[119][120]=0;
index_VN[120][120]=1;
index_VN[120][121]=0;
index_VN[121][121]=1;
index_VN[121][122]=0;
index_VN[122][122]=1;
index_VN[122][123]=0;
index_VN[123][123]=1;
index_VN[123][124]=0;
index_VN[124][124]=1;
index_VN[124][125]=0;
index_VN[125][125]=1;
index_VN[125][126]=0;
index_VN[126][126]=1;
index_VN[126][127]=0;
index_VN[127][127]=1;
index_VN[128][128]=0;
index_VN[255][128]=1;
index_VN[128][129]=0;
index_VN[129][129]=1;
index_VN[129][130]=0;
index_VN[130][130]=1;
index_VN[130][131]=0;
index_VN[131][131]=1;
index_VN[131][132]=0;
index_VN[132][132]=1;
index_VN[132][133]=0;
index_VN[133][133]=1;
index_VN[133][134]=0;
index_VN[134][134]=1;
index_VN[134][135]=0;
index_VN[135][135]=1;
index_VN[135][136]=0;
index_VN[136][136]=1;
index_VN[136][137]=0;
index_VN[137][137]=1;
index_VN[137][138]=0;
index_VN[138][138]=1;
index_VN[138][139]=0;
index_VN[139][139]=1;
index_VN[139][140]=0;
index_VN[140][140]=1;
index_VN[140][141]=0;
index_VN[141][141]=1;
index_VN[141][142]=0;
index_VN[142][142]=1;
index_VN[142][143]=0;
index_VN[143][143]=1;
index_VN[143][144]=0;
index_VN[144][144]=1;
index_VN[144][145]=0;
index_VN[145][145]=1;
index_VN[145][146]=0;
index_VN[146][146]=1;
index_VN[146][147]=0;
index_VN[147][147]=1;
index_VN[147][148]=0;
index_VN[148][148]=1;
index_VN[148][149]=0;
index_VN[149][149]=1;
index_VN[149][150]=0;
index_VN[150][150]=1;
index_VN[150][151]=0;
index_VN[151][151]=1;
index_VN[151][152]=0;
index_VN[152][152]=1;
index_VN[152][153]=0;
index_VN[153][153]=1;
index_VN[153][154]=0;
index_VN[154][154]=1;
index_VN[154][155]=0;
index_VN[155][155]=1;
index_VN[155][156]=0;
index_VN[156][156]=1;
index_VN[156][157]=0;
index_VN[157][157]=1;
index_VN[157][158]=0;
index_VN[158][158]=1;
index_VN[158][159]=0;
index_VN[159][159]=1;
index_VN[159][160]=0;
index_VN[160][160]=1;
index_VN[160][161]=0;
index_VN[161][161]=1;
index_VN[161][162]=0;
index_VN[162][162]=1;
index_VN[162][163]=0;
index_VN[163][163]=1;
index_VN[163][164]=0;
index_VN[164][164]=1;
index_VN[164][165]=0;
index_VN[165][165]=1;
index_VN[165][166]=0;
index_VN[166][166]=1;
index_VN[166][167]=0;
index_VN[167][167]=1;
index_VN[167][168]=0;
index_VN[168][168]=1;
index_VN[168][169]=0;
index_VN[169][169]=1;
index_VN[169][170]=0;
index_VN[170][170]=1;
index_VN[170][171]=0;
index_VN[171][171]=1;
index_VN[171][172]=0;
index_VN[172][172]=1;
index_VN[172][173]=0;
index_VN[173][173]=1;
index_VN[173][174]=0;
index_VN[174][174]=1;
index_VN[174][175]=0;
index_VN[175][175]=1;
index_VN[175][176]=0;
index_VN[176][176]=1;
index_VN[176][177]=0;
index_VN[177][177]=1;
index_VN[177][178]=0;
index_VN[178][178]=1;
index_VN[178][179]=0;
index_VN[179][179]=1;
index_VN[179][180]=0;
index_VN[180][180]=1;
index_VN[180][181]=0;
index_VN[181][181]=1;
index_VN[181][182]=0;
index_VN[182][182]=1;
index_VN[182][183]=0;
index_VN[183][183]=1;
index_VN[183][184]=0;
index_VN[184][184]=1;
index_VN[184][185]=0;
index_VN[185][185]=1;
index_VN[185][186]=0;
index_VN[186][186]=1;
index_VN[186][187]=0;
index_VN[187][187]=1;
index_VN[187][188]=0;
index_VN[188][188]=1;
index_VN[188][189]=0;
index_VN[189][189]=1;
index_VN[189][190]=0;
index_VN[190][190]=1;
index_VN[190][191]=0;
index_VN[191][191]=1;
index_VN[191][192]=0;
index_VN[192][192]=1;
index_VN[192][193]=0;
index_VN[193][193]=1;
index_VN[193][194]=0;
index_VN[194][194]=1;
index_VN[194][195]=0;
index_VN[195][195]=1;
index_VN[195][196]=0;
index_VN[196][196]=1;
index_VN[196][197]=0;
index_VN[197][197]=1;
index_VN[197][198]=0;
index_VN[198][198]=1;
index_VN[198][199]=0;
index_VN[199][199]=1;
index_VN[199][200]=0;
index_VN[200][200]=1;
index_VN[200][201]=0;
index_VN[201][201]=1;
index_VN[201][202]=0;
index_VN[202][202]=1;
index_VN[202][203]=0;
index_VN[203][203]=1;
index_VN[203][204]=0;
index_VN[204][204]=1;
index_VN[204][205]=0;
index_VN[205][205]=1;
index_VN[205][206]=0;
index_VN[206][206]=1;
index_VN[206][207]=0;
index_VN[207][207]=1;
index_VN[207][208]=0;
index_VN[208][208]=1;
index_VN[208][209]=0;
index_VN[209][209]=1;
index_VN[209][210]=0;
index_VN[210][210]=1;
index_VN[210][211]=0;
index_VN[211][211]=1;
index_VN[211][212]=0;
index_VN[212][212]=1;
index_VN[212][213]=0;
index_VN[213][213]=1;
index_VN[213][214]=0;
index_VN[214][214]=1;
index_VN[214][215]=0;
index_VN[215][215]=1;
index_VN[215][216]=0;
index_VN[216][216]=1;
index_VN[216][217]=0;
index_VN[217][217]=1;
index_VN[217][218]=0;
index_VN[218][218]=1;
index_VN[218][219]=0;
index_VN[219][219]=1;
index_VN[219][220]=0;
index_VN[220][220]=1;
index_VN[220][221]=0;
index_VN[221][221]=1;
index_VN[221][222]=0;
index_VN[222][222]=1;
index_VN[222][223]=0;
index_VN[223][223]=1;
index_VN[223][224]=0;
index_VN[224][224]=1;
index_VN[224][225]=0;
index_VN[225][225]=1;
index_VN[225][226]=0;
index_VN[226][226]=1;
index_VN[226][227]=0;
index_VN[227][227]=1;
index_VN[227][228]=0;
index_VN[228][228]=1;
index_VN[228][229]=0;
index_VN[229][229]=1;
index_VN[229][230]=0;
index_VN[230][230]=1;
index_VN[230][231]=0;
index_VN[231][231]=1;
index_VN[231][232]=0;
index_VN[232][232]=1;
index_VN[232][233]=0;
index_VN[233][233]=1;
index_VN[233][234]=0;
index_VN[234][234]=1;
index_VN[234][235]=0;
index_VN[235][235]=1;
index_VN[235][236]=0;
index_VN[236][236]=1;
index_VN[236][237]=0;
index_VN[237][237]=1;
index_VN[237][238]=0;
index_VN[238][238]=1;
index_VN[238][239]=0;
index_VN[239][239]=1;
index_VN[239][240]=0;
index_VN[240][240]=1;
index_VN[240][241]=0;
index_VN[241][241]=1;
index_VN[241][242]=0;
index_VN[242][242]=1;
index_VN[242][243]=0;
index_VN[243][243]=1;
index_VN[243][244]=0;
index_VN[244][244]=1;
index_VN[244][245]=0;
index_VN[245][245]=1;
index_VN[245][246]=0;
index_VN[246][246]=1;
index_VN[246][247]=0;
index_VN[247][247]=1;
index_VN[247][248]=0;
index_VN[248][248]=1;
index_VN[248][249]=0;
index_VN[249][249]=1;
index_VN[249][250]=0;
index_VN[250][250]=1;
index_VN[250][251]=0;
index_VN[251][251]=1;
index_VN[251][252]=0;
index_VN[252][252]=1;
index_VN[252][253]=0;
index_VN[253][253]=1;
index_VN[253][254]=0;
index_VN[254][254]=1;
index_VN[254][255]=0;
index_VN[255][255]=1;
index_VN[0][256]=0;
index_VN[141][256]=1;
index_VN[1][257]=0;
index_VN[132][257]=1;
index_VN[2][258]=0;
index_VN[251][258]=1;
index_VN[3][259]=0;
index_VN[148][259]=1;
index_VN[4][260]=0;
index_VN[243][260]=1;
index_VN[5][261]=0;
index_VN[156][261]=1;
index_VN[6][262]=0;
index_VN[165][262]=1;
index_VN[7][263]=0;
index_VN[236][263]=1;
index_VN[8][264]=0;
index_VN[135][264]=1;
index_VN[9][265]=0;
index_VN[172][265]=1;
index_VN[10][266]=0;
index_VN[145][266]=1;
index_VN[11][267]=0;
index_VN[246][267]=1;
index_VN[12][268]=0;
index_VN[129][268]=1;
index_VN[13][269]=0;
index_VN[152][269]=1;
index_VN[14][270]=0;
index_VN[177][270]=1;
index_VN[15][271]=0;
index_VN[238][271]=1;
index_VN[16][272]=0;
index_VN[159][272]=1;
index_VN[17][273]=0;
index_VN[184][273]=1;
index_VN[18][274]=0;
index_VN[231][274]=1;
index_VN[19][275]=0;
index_VN[254][275]=1;
index_VN[20][276]=0;
index_VN[223][276]=1;
index_VN[21][277]=0;
index_VN[142][277]=1;
index_VN[22][278]=0;
index_VN[153][278]=1;
index_VN[23][279]=0;
index_VN[170][279]=1;
index_VN[24][280]=0;
index_VN[187][280]=1;
index_VN[25][281]=0;
index_VN[242][281]=1;
index_VN[26][282]=0;
index_VN[195][282]=1;
index_VN[27][283]=0;
index_VN[230][283]=1;
index_VN[28][284]=0;
index_VN[219][284]=1;
index_VN[29][285]=0;
index_VN[174][285]=1;
index_VN[30][286]=0;
index_VN[211][286]=1;
index_VN[31][287]=0;
index_VN[200][287]=1;
index_VN[32][288]=0;
index_VN[167][288]=1;
index_VN[33][289]=0;
index_VN[138][289]=1;
index_VN[34][290]=0;
index_VN[247][290]=1;
index_VN[35][291]=0;
index_VN[228][291]=1;
index_VN[36][292]=0;
index_VN[189][292]=1;
index_VN[37][293]=0;
index_VN[150][293]=1;
index_VN[38][294]=0;
index_VN[163][294]=1;
index_VN[39][295]=0;
index_VN[198][295]=1;
index_VN[40][296]=0;
index_VN[217][296]=1;
index_VN[41][297]=0;
index_VN[134][297]=1;
index_VN[42][298]=0;
index_VN[209][298]=1;
index_VN[43][299]=0;
index_VN[186][299]=1;
index_VN[44][300]=0;
index_VN[147][300]=1;
index_VN[45][301]=0;
index_VN[224][301]=1;
index_VN[46][302]=0;
index_VN[175][302]=1;
index_VN[47][303]=0;
index_VN[248][303]=1;
index_VN[48][304]=0;
index_VN[205][304]=1;
index_VN[49][305]=0;
index_VN[158][305]=1;
index_VN[50][306]=0;
index_VN[197][306]=1;
index_VN[51][307]=0;
index_VN[144][307]=1;
index_VN[52][308]=0;
index_VN[181][308]=1;
index_VN[53][309]=0;
index_VN[214][309]=1;
index_VN[54][310]=0;
index_VN[239][310]=1;
index_VN[55][311]=0;
index_VN[190][311]=1;
index_VN[56][312]=0;
index_VN[253][312]=1;
index_VN[57][313]=0;
index_VN[208][313]=1;
index_VN[58][314]=0;
index_VN[139][314]=1;
index_VN[59][315]=0;
index_VN[162][315]=1;
index_VN[60][316]=0;
index_VN[225][316]=1;
index_VN[61][317]=0;
index_VN[244][317]=1;
index_VN[62][318]=0;
index_VN[203][318]=1;
index_VN[63][319]=0;
index_VN[178][319]=1;
index_VN[64][320]=0;
index_VN[133][320]=1;
index_VN[65][321]=0;
index_VN[194][321]=1;
index_VN[66][322]=0;
index_VN[155][322]=1;
index_VN[67][323]=0;
index_VN[212][323]=1;
index_VN[68][324]=0;
index_VN[255][324]=1;
index_VN[69][325]=0;
index_VN[149][325]=1;
index_VN[70][326]=0;
index_VN[136][326]=1;
index_VN[71][327]=0;
index_VN[183][327]=1;
index_VN[72][328]=0;
index_VN[221][328]=1;
index_VN[73][329]=0;
index_VN[250][329]=1;
index_VN[74][330]=0;
index_VN[168][330]=1;
index_VN[75][331]=0;
index_VN[215][331]=1;
index_VN[76][332]=0;
index_VN[226][332]=1;
index_VN[77][333]=0;
index_VN[234][333]=1;
index_VN[78][334]=0;
index_VN[128][334]=1;
index_VN[79][335]=0;
index_VN[196][335]=1;
index_VN[80][336]=0;
index_VN[140][336]=1;
index_VN[81][337]=0;
index_VN[173][337]=1;
index_VN[82][338]=0;
index_VN[182][338]=1;
index_VN[83][339]=0;
index_VN[154][339]=1;
index_VN[84][340]=0;
index_VN[202][340]=1;
index_VN[85][341]=0;
index_VN[191][341]=1;
index_VN[86][342]=0;
index_VN[131][342]=1;
index_VN[87][343]=0;
index_VN[169][343]=1;
index_VN[88][344]=0;
index_VN[161][344]=1;
index_VN[89][345]=0;
index_VN[180][345]=1;
index_VN[90][346]=0;
index_VN[232][346]=1;
index_VN[91][347]=0;
index_VN[245][347]=1;
index_VN[92][348]=0;
index_VN[216][348]=1;
index_VN[93][349]=0;
index_VN[192][349]=1;
index_VN[94][350]=0;
index_VN[143][350]=1;
index_VN[95][351]=0;
index_VN[164][351]=1;
index_VN[96][352]=0;
index_VN[252][352]=1;
index_VN[97][353]=0;
index_VN[176][353]=1;
index_VN[98][354]=0;
index_VN[233][354]=1;
index_VN[99][355]=0;
index_VN[137][355]=1;
index_VN[100][356]=0;
index_VN[157][356]=1;
index_VN[101][357]=0;
index_VN[188][357]=1;
index_VN[102][358]=0;
index_VN[220][358]=1;
index_VN[103][359]=0;
index_VN[130][359]=1;
index_VN[104][360]=0;
index_VN[206][360]=1;
index_VN[105][361]=0;
index_VN[237][361]=1;
index_VN[106][362]=0;
index_VN[229][362]=1;
index_VN[107][363]=0;
index_VN[146][363]=1;
index_VN[108][364]=0;
index_VN[201][364]=1;
index_VN[109][365]=0;
index_VN[249][365]=1;
index_VN[110][366]=0;
index_VN[241][366]=1;
index_VN[111][367]=0;
index_VN[151][367]=1;
index_VN[112][368]=0;
index_VN[210][368]=1;
index_VN[113][369]=0;
index_VN[235][369]=1;
index_VN[114][370]=0;
index_VN[193][370]=1;
index_VN[115][371]=0;
index_VN[160][371]=1;
index_VN[116][372]=0;
index_VN[222][372]=1;
index_VN[117][373]=0;
index_VN[199][373]=1;
index_VN[118][374]=0;
index_VN[171][374]=1;
index_VN[119][375]=0;
index_VN[207][375]=1;
index_VN[120][376]=0;
index_VN[179][376]=1;
index_VN[121][377]=0;
index_VN[218][377]=1;
index_VN[122][378]=0;
index_VN[166][378]=1;
index_VN[123][379]=0;
index_VN[240][379]=1;
index_VN[124][380]=0;
index_VN[227][380]=1;
index_VN[125][381]=0;
index_VN[185][381]=1;
index_VN[126][382]=0;
index_VN[204][382]=1;
index_VN[127][383]=0;
index_VN[213][383]=1;

/* MAGICS DECLARATIONS*/
index_CN[0][0]=0;
index_CN[0][1]=1;
index_CN[0][256]=2;
index_CN[1][1]=0;
index_CN[1][2]=1;
index_CN[1][257]=2;
index_CN[2][2]=0;
index_CN[2][3]=1;
index_CN[2][258]=2;
index_CN[3][3]=0;
index_CN[3][4]=1;
index_CN[3][259]=2;
index_CN[4][4]=0;
index_CN[4][5]=1;
index_CN[4][260]=2;
index_CN[5][5]=0;
index_CN[5][6]=1;
index_CN[5][261]=2;
index_CN[6][6]=0;
index_CN[6][7]=1;
index_CN[6][262]=2;
index_CN[7][7]=0;
index_CN[7][8]=1;
index_CN[7][263]=2;
index_CN[8][8]=0;
index_CN[8][9]=1;
index_CN[8][264]=2;
index_CN[9][9]=0;
index_CN[9][10]=1;
index_CN[9][265]=2;
index_CN[10][10]=0;
index_CN[10][11]=1;
index_CN[10][266]=2;
index_CN[11][11]=0;
index_CN[11][12]=1;
index_CN[11][267]=2;
index_CN[12][12]=0;
index_CN[12][13]=1;
index_CN[12][268]=2;
index_CN[13][13]=0;
index_CN[13][14]=1;
index_CN[13][269]=2;
index_CN[14][14]=0;
index_CN[14][15]=1;
index_CN[14][270]=2;
index_CN[15][15]=0;
index_CN[15][16]=1;
index_CN[15][271]=2;
index_CN[16][16]=0;
index_CN[16][17]=1;
index_CN[16][272]=2;
index_CN[17][17]=0;
index_CN[17][18]=1;
index_CN[17][273]=2;
index_CN[18][18]=0;
index_CN[18][19]=1;
index_CN[18][274]=2;
index_CN[19][19]=0;
index_CN[19][20]=1;
index_CN[19][275]=2;
index_CN[20][20]=0;
index_CN[20][21]=1;
index_CN[20][276]=2;
index_CN[21][21]=0;
index_CN[21][22]=1;
index_CN[21][277]=2;
index_CN[22][22]=0;
index_CN[22][23]=1;
index_CN[22][278]=2;
index_CN[23][23]=0;
index_CN[23][24]=1;
index_CN[23][279]=2;
index_CN[24][24]=0;
index_CN[24][25]=1;
index_CN[24][280]=2;
index_CN[25][25]=0;
index_CN[25][26]=1;
index_CN[25][281]=2;
index_CN[26][26]=0;
index_CN[26][27]=1;
index_CN[26][282]=2;
index_CN[27][27]=0;
index_CN[27][28]=1;
index_CN[27][283]=2;
index_CN[28][28]=0;
index_CN[28][29]=1;
index_CN[28][284]=2;
index_CN[29][29]=0;
index_CN[29][30]=1;
index_CN[29][285]=2;
index_CN[30][30]=0;
index_CN[30][31]=1;
index_CN[30][286]=2;
index_CN[31][31]=0;
index_CN[31][32]=1;
index_CN[31][287]=2;
index_CN[32][32]=0;
index_CN[32][33]=1;
index_CN[32][288]=2;
index_CN[33][33]=0;
index_CN[33][34]=1;
index_CN[33][289]=2;
index_CN[34][34]=0;
index_CN[34][35]=1;
index_CN[34][290]=2;
index_CN[35][35]=0;
index_CN[35][36]=1;
index_CN[35][291]=2;
index_CN[36][36]=0;
index_CN[36][37]=1;
index_CN[36][292]=2;
index_CN[37][37]=0;
index_CN[37][38]=1;
index_CN[37][293]=2;
index_CN[38][38]=0;
index_CN[38][39]=1;
index_CN[38][294]=2;
index_CN[39][39]=0;
index_CN[39][40]=1;
index_CN[39][295]=2;
index_CN[40][40]=0;
index_CN[40][41]=1;
index_CN[40][296]=2;
index_CN[41][41]=0;
index_CN[41][42]=1;
index_CN[41][297]=2;
index_CN[42][42]=0;
index_CN[42][43]=1;
index_CN[42][298]=2;
index_CN[43][43]=0;
index_CN[43][44]=1;
index_CN[43][299]=2;
index_CN[44][44]=0;
index_CN[44][45]=1;
index_CN[44][300]=2;
index_CN[45][45]=0;
index_CN[45][46]=1;
index_CN[45][301]=2;
index_CN[46][46]=0;
index_CN[46][47]=1;
index_CN[46][302]=2;
index_CN[47][47]=0;
index_CN[47][48]=1;
index_CN[47][303]=2;
index_CN[48][48]=0;
index_CN[48][49]=1;
index_CN[48][304]=2;
index_CN[49][49]=0;
index_CN[49][50]=1;
index_CN[49][305]=2;
index_CN[50][50]=0;
index_CN[50][51]=1;
index_CN[50][306]=2;
index_CN[51][51]=0;
index_CN[51][52]=1;
index_CN[51][307]=2;
index_CN[52][52]=0;
index_CN[52][53]=1;
index_CN[52][308]=2;
index_CN[53][53]=0;
index_CN[53][54]=1;
index_CN[53][309]=2;
index_CN[54][54]=0;
index_CN[54][55]=1;
index_CN[54][310]=2;
index_CN[55][55]=0;
index_CN[55][56]=1;
index_CN[55][311]=2;
index_CN[56][56]=0;
index_CN[56][57]=1;
index_CN[56][312]=2;
index_CN[57][57]=0;
index_CN[57][58]=1;
index_CN[57][313]=2;
index_CN[58][58]=0;
index_CN[58][59]=1;
index_CN[58][314]=2;
index_CN[59][59]=0;
index_CN[59][60]=1;
index_CN[59][315]=2;
index_CN[60][60]=0;
index_CN[60][61]=1;
index_CN[60][316]=2;
index_CN[61][61]=0;
index_CN[61][62]=1;
index_CN[61][317]=2;
index_CN[62][62]=0;
index_CN[62][63]=1;
index_CN[62][318]=2;
index_CN[63][63]=0;
index_CN[63][64]=1;
index_CN[63][319]=2;
index_CN[64][64]=0;
index_CN[64][65]=1;
index_CN[64][320]=2;
index_CN[65][65]=0;
index_CN[65][66]=1;
index_CN[65][321]=2;
index_CN[66][66]=0;
index_CN[66][67]=1;
index_CN[66][322]=2;
index_CN[67][67]=0;
index_CN[67][68]=1;
index_CN[67][323]=2;
index_CN[68][68]=0;
index_CN[68][69]=1;
index_CN[68][324]=2;
index_CN[69][69]=0;
index_CN[69][70]=1;
index_CN[69][325]=2;
index_CN[70][70]=0;
index_CN[70][71]=1;
index_CN[70][326]=2;
index_CN[71][71]=0;
index_CN[71][72]=1;
index_CN[71][327]=2;
index_CN[72][72]=0;
index_CN[72][73]=1;
index_CN[72][328]=2;
index_CN[73][73]=0;
index_CN[73][74]=1;
index_CN[73][329]=2;
index_CN[74][74]=0;
index_CN[74][75]=1;
index_CN[74][330]=2;
index_CN[75][75]=0;
index_CN[75][76]=1;
index_CN[75][331]=2;
index_CN[76][76]=0;
index_CN[76][77]=1;
index_CN[76][332]=2;
index_CN[77][77]=0;
index_CN[77][78]=1;
index_CN[77][333]=2;
index_CN[78][78]=0;
index_CN[78][79]=1;
index_CN[78][334]=2;
index_CN[79][79]=0;
index_CN[79][80]=1;
index_CN[79][335]=2;
index_CN[80][80]=0;
index_CN[80][81]=1;
index_CN[80][336]=2;
index_CN[81][81]=0;
index_CN[81][82]=1;
index_CN[81][337]=2;
index_CN[82][82]=0;
index_CN[82][83]=1;
index_CN[82][338]=2;
index_CN[83][83]=0;
index_CN[83][84]=1;
index_CN[83][339]=2;
index_CN[84][84]=0;
index_CN[84][85]=1;
index_CN[84][340]=2;
index_CN[85][85]=0;
index_CN[85][86]=1;
index_CN[85][341]=2;
index_CN[86][86]=0;
index_CN[86][87]=1;
index_CN[86][342]=2;
index_CN[87][87]=0;
index_CN[87][88]=1;
index_CN[87][343]=2;
index_CN[88][88]=0;
index_CN[88][89]=1;
index_CN[88][344]=2;
index_CN[89][89]=0;
index_CN[89][90]=1;
index_CN[89][345]=2;
index_CN[90][90]=0;
index_CN[90][91]=1;
index_CN[90][346]=2;
index_CN[91][91]=0;
index_CN[91][92]=1;
index_CN[91][347]=2;
index_CN[92][92]=0;
index_CN[92][93]=1;
index_CN[92][348]=2;
index_CN[93][93]=0;
index_CN[93][94]=1;
index_CN[93][349]=2;
index_CN[94][94]=0;
index_CN[94][95]=1;
index_CN[94][350]=2;
index_CN[95][95]=0;
index_CN[95][96]=1;
index_CN[95][351]=2;
index_CN[96][96]=0;
index_CN[96][97]=1;
index_CN[96][352]=2;
index_CN[97][97]=0;
index_CN[97][98]=1;
index_CN[97][353]=2;
index_CN[98][98]=0;
index_CN[98][99]=1;
index_CN[98][354]=2;
index_CN[99][99]=0;
index_CN[99][100]=1;
index_CN[99][355]=2;
index_CN[100][100]=0;
index_CN[100][101]=1;
index_CN[100][356]=2;
index_CN[101][101]=0;
index_CN[101][102]=1;
index_CN[101][357]=2;
index_CN[102][102]=0;
index_CN[102][103]=1;
index_CN[102][358]=2;
index_CN[103][103]=0;
index_CN[103][104]=1;
index_CN[103][359]=2;
index_CN[104][104]=0;
index_CN[104][105]=1;
index_CN[104][360]=2;
index_CN[105][105]=0;
index_CN[105][106]=1;
index_CN[105][361]=2;
index_CN[106][106]=0;
index_CN[106][107]=1;
index_CN[106][362]=2;
index_CN[107][107]=0;
index_CN[107][108]=1;
index_CN[107][363]=2;
index_CN[108][108]=0;
index_CN[108][109]=1;
index_CN[108][364]=2;
index_CN[109][109]=0;
index_CN[109][110]=1;
index_CN[109][365]=2;
index_CN[110][110]=0;
index_CN[110][111]=1;
index_CN[110][366]=2;
index_CN[111][111]=0;
index_CN[111][112]=1;
index_CN[111][367]=2;
index_CN[112][112]=0;
index_CN[112][113]=1;
index_CN[112][368]=2;
index_CN[113][113]=0;
index_CN[113][114]=1;
index_CN[113][369]=2;
index_CN[114][114]=0;
index_CN[114][115]=1;
index_CN[114][370]=2;
index_CN[115][115]=0;
index_CN[115][116]=1;
index_CN[115][371]=2;
index_CN[116][116]=0;
index_CN[116][117]=1;
index_CN[116][372]=2;
index_CN[117][117]=0;
index_CN[117][118]=1;
index_CN[117][373]=2;
index_CN[118][118]=0;
index_CN[118][119]=1;
index_CN[118][374]=2;
index_CN[119][119]=0;
index_CN[119][120]=1;
index_CN[119][375]=2;
index_CN[120][120]=0;
index_CN[120][121]=1;
index_CN[120][376]=2;
index_CN[121][121]=0;
index_CN[121][122]=1;
index_CN[121][377]=2;
index_CN[122][122]=0;
index_CN[122][123]=1;
index_CN[122][378]=2;
index_CN[123][123]=0;
index_CN[123][124]=1;
index_CN[123][379]=2;
index_CN[124][124]=0;
index_CN[124][125]=1;
index_CN[124][380]=2;
index_CN[125][125]=0;
index_CN[125][126]=1;
index_CN[125][381]=2;
index_CN[126][126]=0;
index_CN[126][127]=1;
index_CN[126][382]=2;
index_CN[127][0]=0;
index_CN[127][127]=1;
index_CN[127][383]=2;
index_CN[128][128]=0;
index_CN[128][129]=1;
index_CN[128][334]=2;
index_CN[129][129]=0;
index_CN[129][130]=1;
index_CN[129][268]=2;
index_CN[130][130]=0;
index_CN[130][131]=1;
index_CN[130][359]=2;
index_CN[131][131]=0;
index_CN[131][132]=1;
index_CN[131][342]=2;
index_CN[132][132]=0;
index_CN[132][133]=1;
index_CN[132][257]=2;
index_CN[133][133]=0;
index_CN[133][134]=1;
index_CN[133][320]=2;
index_CN[134][134]=0;
index_CN[134][135]=1;
index_CN[134][297]=2;
index_CN[135][135]=0;
index_CN[135][136]=1;
index_CN[135][264]=2;
index_CN[136][136]=0;
index_CN[136][137]=1;
index_CN[136][326]=2;
index_CN[137][137]=0;
index_CN[137][138]=1;
index_CN[137][355]=2;
index_CN[138][138]=0;
index_CN[138][139]=1;
index_CN[138][289]=2;
index_CN[139][139]=0;
index_CN[139][140]=1;
index_CN[139][314]=2;
index_CN[140][140]=0;
index_CN[140][141]=1;
index_CN[140][336]=2;
index_CN[141][141]=0;
index_CN[141][142]=1;
index_CN[141][256]=2;
index_CN[142][142]=0;
index_CN[142][143]=1;
index_CN[142][277]=2;
index_CN[143][143]=0;
index_CN[143][144]=1;
index_CN[143][350]=2;
index_CN[144][144]=0;
index_CN[144][145]=1;
index_CN[144][307]=2;
index_CN[145][145]=0;
index_CN[145][146]=1;
index_CN[145][266]=2;
index_CN[146][146]=0;
index_CN[146][147]=1;
index_CN[146][363]=2;
index_CN[147][147]=0;
index_CN[147][148]=1;
index_CN[147][300]=2;
index_CN[148][148]=0;
index_CN[148][149]=1;
index_CN[148][259]=2;
index_CN[149][149]=0;
index_CN[149][150]=1;
index_CN[149][325]=2;
index_CN[150][150]=0;
index_CN[150][151]=1;
index_CN[150][293]=2;
index_CN[151][151]=0;
index_CN[151][152]=1;
index_CN[151][367]=2;
index_CN[152][152]=0;
index_CN[152][153]=1;
index_CN[152][269]=2;
index_CN[153][153]=0;
index_CN[153][154]=1;
index_CN[153][278]=2;
index_CN[154][154]=0;
index_CN[154][155]=1;
index_CN[154][339]=2;
index_CN[155][155]=0;
index_CN[155][156]=1;
index_CN[155][322]=2;
index_CN[156][156]=0;
index_CN[156][157]=1;
index_CN[156][261]=2;
index_CN[157][157]=0;
index_CN[157][158]=1;
index_CN[157][356]=2;
index_CN[158][158]=0;
index_CN[158][159]=1;
index_CN[158][305]=2;
index_CN[159][159]=0;
index_CN[159][160]=1;
index_CN[159][272]=2;
index_CN[160][160]=0;
index_CN[160][161]=1;
index_CN[160][371]=2;
index_CN[161][161]=0;
index_CN[161][162]=1;
index_CN[161][344]=2;
index_CN[162][162]=0;
index_CN[162][163]=1;
index_CN[162][315]=2;
index_CN[163][163]=0;
index_CN[163][164]=1;
index_CN[163][294]=2;
index_CN[164][164]=0;
index_CN[164][165]=1;
index_CN[164][351]=2;
index_CN[165][165]=0;
index_CN[165][166]=1;
index_CN[165][262]=2;
index_CN[166][166]=0;
index_CN[166][167]=1;
index_CN[166][378]=2;
index_CN[167][167]=0;
index_CN[167][168]=1;
index_CN[167][288]=2;
index_CN[168][168]=0;
index_CN[168][169]=1;
index_CN[168][330]=2;
index_CN[169][169]=0;
index_CN[169][170]=1;
index_CN[169][343]=2;
index_CN[170][170]=0;
index_CN[170][171]=1;
index_CN[170][279]=2;
index_CN[171][171]=0;
index_CN[171][172]=1;
index_CN[171][374]=2;
index_CN[172][172]=0;
index_CN[172][173]=1;
index_CN[172][265]=2;
index_CN[173][173]=0;
index_CN[173][174]=1;
index_CN[173][337]=2;
index_CN[174][174]=0;
index_CN[174][175]=1;
index_CN[174][285]=2;
index_CN[175][175]=0;
index_CN[175][176]=1;
index_CN[175][302]=2;
index_CN[176][176]=0;
index_CN[176][177]=1;
index_CN[176][353]=2;
index_CN[177][177]=0;
index_CN[177][178]=1;
index_CN[177][270]=2;
index_CN[178][178]=0;
index_CN[178][179]=1;
index_CN[178][319]=2;
index_CN[179][179]=0;
index_CN[179][180]=1;
index_CN[179][376]=2;
index_CN[180][180]=0;
index_CN[180][181]=1;
index_CN[180][345]=2;
index_CN[181][181]=0;
index_CN[181][182]=1;
index_CN[181][308]=2;
index_CN[182][182]=0;
index_CN[182][183]=1;
index_CN[182][338]=2;
index_CN[183][183]=0;
index_CN[183][184]=1;
index_CN[183][327]=2;
index_CN[184][184]=0;
index_CN[184][185]=1;
index_CN[184][273]=2;
index_CN[185][185]=0;
index_CN[185][186]=1;
index_CN[185][381]=2;
index_CN[186][186]=0;
index_CN[186][187]=1;
index_CN[186][299]=2;
index_CN[187][187]=0;
index_CN[187][188]=1;
index_CN[187][280]=2;
index_CN[188][188]=0;
index_CN[188][189]=1;
index_CN[188][357]=2;
index_CN[189][189]=0;
index_CN[189][190]=1;
index_CN[189][292]=2;
index_CN[190][190]=0;
index_CN[190][191]=1;
index_CN[190][311]=2;
index_CN[191][191]=0;
index_CN[191][192]=1;
index_CN[191][341]=2;
index_CN[192][192]=0;
index_CN[192][193]=1;
index_CN[192][349]=2;
index_CN[193][193]=0;
index_CN[193][194]=1;
index_CN[193][370]=2;
index_CN[194][194]=0;
index_CN[194][195]=1;
index_CN[194][321]=2;
index_CN[195][195]=0;
index_CN[195][196]=1;
index_CN[195][282]=2;
index_CN[196][196]=0;
index_CN[196][197]=1;
index_CN[196][335]=2;
index_CN[197][197]=0;
index_CN[197][198]=1;
index_CN[197][306]=2;
index_CN[198][198]=0;
index_CN[198][199]=1;
index_CN[198][295]=2;
index_CN[199][199]=0;
index_CN[199][200]=1;
index_CN[199][373]=2;
index_CN[200][200]=0;
index_CN[200][201]=1;
index_CN[200][287]=2;
index_CN[201][201]=0;
index_CN[201][202]=1;
index_CN[201][364]=2;
index_CN[202][202]=0;
index_CN[202][203]=1;
index_CN[202][340]=2;
index_CN[203][203]=0;
index_CN[203][204]=1;
index_CN[203][318]=2;
index_CN[204][204]=0;
index_CN[204][205]=1;
index_CN[204][382]=2;
index_CN[205][205]=0;
index_CN[205][206]=1;
index_CN[205][304]=2;
index_CN[206][206]=0;
index_CN[206][207]=1;
index_CN[206][360]=2;
index_CN[207][207]=0;
index_CN[207][208]=1;
index_CN[207][375]=2;
index_CN[208][208]=0;
index_CN[208][209]=1;
index_CN[208][313]=2;
index_CN[209][209]=0;
index_CN[209][210]=1;
index_CN[209][298]=2;
index_CN[210][210]=0;
index_CN[210][211]=1;
index_CN[210][368]=2;
index_CN[211][211]=0;
index_CN[211][212]=1;
index_CN[211][286]=2;
index_CN[212][212]=0;
index_CN[212][213]=1;
index_CN[212][323]=2;
index_CN[213][213]=0;
index_CN[213][214]=1;
index_CN[213][383]=2;
index_CN[214][214]=0;
index_CN[214][215]=1;
index_CN[214][309]=2;
index_CN[215][215]=0;
index_CN[215][216]=1;
index_CN[215][331]=2;
index_CN[216][216]=0;
index_CN[216][217]=1;
index_CN[216][348]=2;
index_CN[217][217]=0;
index_CN[217][218]=1;
index_CN[217][296]=2;
index_CN[218][218]=0;
index_CN[218][219]=1;
index_CN[218][377]=2;
index_CN[219][219]=0;
index_CN[219][220]=1;
index_CN[219][284]=2;
index_CN[220][220]=0;
index_CN[220][221]=1;
index_CN[220][358]=2;
index_CN[221][221]=0;
index_CN[221][222]=1;
index_CN[221][328]=2;
index_CN[222][222]=0;
index_CN[222][223]=1;
index_CN[222][372]=2;
index_CN[223][223]=0;
index_CN[223][224]=1;
index_CN[223][276]=2;
index_CN[224][224]=0;
index_CN[224][225]=1;
index_CN[224][301]=2;
index_CN[225][225]=0;
index_CN[225][226]=1;
index_CN[225][316]=2;
index_CN[226][226]=0;
index_CN[226][227]=1;
index_CN[226][332]=2;
index_CN[227][227]=0;
index_CN[227][228]=1;
index_CN[227][380]=2;
index_CN[228][228]=0;
index_CN[228][229]=1;
index_CN[228][291]=2;
index_CN[229][229]=0;
index_CN[229][230]=1;
index_CN[229][362]=2;
index_CN[230][230]=0;
index_CN[230][231]=1;
index_CN[230][283]=2;
index_CN[231][231]=0;
index_CN[231][232]=1;
index_CN[231][274]=2;
index_CN[232][232]=0;
index_CN[232][233]=1;
index_CN[232][346]=2;
index_CN[233][233]=0;
index_CN[233][234]=1;
index_CN[233][354]=2;
index_CN[234][234]=0;
index_CN[234][235]=1;
index_CN[234][333]=2;
index_CN[235][235]=0;
index_CN[235][236]=1;
index_CN[235][369]=2;
index_CN[236][236]=0;
index_CN[236][237]=1;
index_CN[236][263]=2;
index_CN[237][237]=0;
index_CN[237][238]=1;
index_CN[237][361]=2;
index_CN[238][238]=0;
index_CN[238][239]=1;
index_CN[238][271]=2;
index_CN[239][239]=0;
index_CN[239][240]=1;
index_CN[239][310]=2;
index_CN[240][240]=0;
index_CN[240][241]=1;
index_CN[240][379]=2;
index_CN[241][241]=0;
index_CN[241][242]=1;
index_CN[241][366]=2;
index_CN[242][242]=0;
index_CN[242][243]=1;
index_CN[242][281]=2;
index_CN[243][243]=0;
index_CN[243][244]=1;
index_CN[243][260]=2;
index_CN[244][244]=0;
index_CN[244][245]=1;
index_CN[244][317]=2;
index_CN[245][245]=0;
index_CN[245][246]=1;
index_CN[245][347]=2;
index_CN[246][246]=0;
index_CN[246][247]=1;
index_CN[246][267]=2;
index_CN[247][247]=0;
index_CN[247][248]=1;
index_CN[247][290]=2;
index_CN[248][248]=0;
index_CN[248][249]=1;
index_CN[248][303]=2;
index_CN[249][249]=0;
index_CN[249][250]=1;
index_CN[249][365]=2;
index_CN[250][250]=0;
index_CN[250][251]=1;
index_CN[250][329]=2;
index_CN[251][251]=0;
index_CN[251][252]=1;
index_CN[251][258]=2;
index_CN[252][252]=0;
index_CN[252][253]=1;
index_CN[252][352]=2;
index_CN[253][253]=0;
index_CN[253][254]=1;
index_CN[253][312]=2;
index_CN[254][254]=0;
index_CN[254][255]=1;
index_CN[254][275]=2;
index_CN[255][128]=0;
index_CN[255][255]=1;
index_CN[255][324]=2;


/* OTHER INITIALIZATIONS*/
row=0;
col=0;
end


else begin
case(state)

`gammaIn: begin
Gamma[row][col]=gamma;

//case(col)
//9'd384: begin

//end
case(row)
QQ: begin
case(col)
9'd383: begin
   state=`alpha_Init;
   c=0;
   a=0;
   col=0;
   end
default: begin
   col=col+1;
   row=0;
end
 endcase
end
default: begin
row=row+1;
end
endcase

                                            



end

/* END OF THE STATE*/


`alpha_Init: begin



     for(c=0;c<2;c=c+1) begin//this is to access row col 
        for(col=0;col<384;col=col+1)// each column is filled
           begin
                row=row_col[c][col];// rowcol is necessary to access only non zero rows of the alpha
                expanded_address=index_VN[row][col];
                 address_index=expanded_address+(col*2);
                 addrAW[address_index]=a;
                 dinA[address_index]=Gamma[a][col];
                 weA[address_index]=1;
               
           end
           
end
case(a)
QQ: begin
 state=`processing_statex;
 a=0;
 end
default: begin
a=a+1;
end
endcase
end


`processing_statex: begin
for(address_index1=0;address_index1<768;address_index1=address_index1+1)
 begin
 weA[address_index1]=0;
 end
for(row=0;row<256;row=row+1)
begin
//col=col_row[row][0];

col=col_row[row][0];
inv_gf(H[row][col],inv_val);
mul_gf(inv_val,0,mul_val);



expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=mul_val;
end

state=`processing_state;
end
`processing_state: begin

for(address_index1=0;address_index1<768;address_index1=address_index1+1)
 begin
 weA[address_index1]=0;
 end
for(row=0;row<256;row=row+1)
begin
col=col_row[row][0];


inv_gf(H[row][col],inv_val);
mul_gf(inv_val,1,mul_val);

expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=mul_val;
end
a=2;
b=0;
state=`F_init1;
end
`F_init1:begin
for(address_index1=0;address_index1<768;address_index1=address_index1+1)
 begin
 weA[address_index1]=0;
 end
for(row=0;row<256;row=row+1)
begin
col=col_row[row][0];
inv_gf(H[row][col],inv_val);
mul_gf(inv_val,a,mul_val);
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=mul_val;
end
for(row=0;row<256;row=row+1)
begin
col=col_row[row][0];
expanded_address=index_VN[row][col];
address_index2=(col*2)+expanded_address;

F[b][0][row]=doutA[address_index2];
end

case(b)
QQ: begin
state=`processing_state1;
for(address_index1=0;address_index1<768;address_index1=address_index1+1)
 begin
 weA[address_index1]=0;
 end
for(row=0;row<256;row=row+1)
begin
col=col_row[row][2];
inv_gf(H[row][col],inv_val);
mul_gf(inv_val,0,mul_val);
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=mul_val;

end

end 
default: begin
b=b+1;
a=a+1;
end
endcase

end



////////

`processing_state1: begin

for(address_index1=0;address_index1<768;address_index1=address_index1+1)
 begin
 weA[address_index1]=0;
 end
for(row=0;row<256;row=row+1)
begin
col=col_row[row][2];
inv_gf(H[row][col],inv_val);
mul_gf(inv_val,1,mul_val);
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=mul_val;
end
a=2;
b=0;


state=`B_init1;
end





`B_init1: begin

for(address_index1=0;address_index1<768;address_index1=address_index1+1)
 begin
 weA[address_index1]=0;
 end
for(row=0;row<256;row=row+1)
begin
col=col_row[row][2];
expanded_address=index_VN[row][col];
inv_gf(H[row][col],inv_val);
mul_gf(inv_val,a,mul_val);
address_index=(col*2)+expanded_address;
addrAR[address_index]=mul_val;
end

for(row=0;row<256;row=row+1)
begin
col=col_row[row][2];

expanded_address=index_VN[row][col];
address_index2=(col*2)+expanded_address;

B[b][2][row]=doutA[address_index2];
end
case(b)
QQ: begin
 state=`processing_state2;
 s=1;
 a=0;
 end
default: begin
b=b+1;
a=a+1;
end
endcase

end

`processing_state2: begin
for(row=0;row<256;row=row+1)
begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=0;
weA[address_index]=0;
end
state=`processing_state3;
end
`processing_state3: begin
for(row=0;row<256;row=row+1)
begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=1;
weA[address_index]=0;
end
a=2;
b=0;
state=`Alphadecide;
end
`Alphadecide: begin
for(row=0;row<256;row=row+1)
begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=a;
weA[address_index]=0;
end

for(row=0;row<256;row=row+1)
begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
AlphaSet[b][row]=doutA[address_index];
end
case(b)
QQ:state=`F_init2;
default:begin
a=a+1;
b=b+1;
end
endcase
end
`F_init2: begin
for(row=0;row<256;row=row+1)begin
col=col_row[row][s];
for(c = 0; c < (QQ+1); c=c+1)begin


						min_F[row][c] = max(F[c][s-1][row],AlphaSet[0][row]);

						for(b = 1; b < (QQ+1); b=b+1)begin
							mul_gf(H[row][col],b,mul_val);
                             add_gf(c,mul_val,a);


							max_F[row][c] = max(F[a][s-1][row], AlphaSet[b][row]);
							min_F[row][c] = min(min_F[row][c], max_F[row][c]);

						end
	//					F[c][s][row] = min_F[row];


					end


end
state=`F_init21;
end
`F_init21: begin

for(row=0;row<256;row=row+1) begin
for(c=0;c<(QQ+1);c=c+1) begin
F[c][s][row]=min_F[row][c];
end

end

case(s)
2:begin
state=`processing_state4;
s=1;
end
default:begin
s=s+1;
state=`processing_state2;
end
endcase
end

`processing_state4: begin
//col=col_row[row][s];
for(row=0;row<256;row=row+1) begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=0;
weA[address_index]=0;
end
state=`processing_state5;
end
`processing_state5: begin
for(row=0;row<256;row=row+1) begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=1;
weA[address_index]=0;
a=2;
b=0;
end
state=`Alphadecide1;
end
`Alphadecide1: begin
for(row=0;row<256;row=row+1)
begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
addrAR[address_index]=a;
weA[address_index]=0;
end

for(row=0;row<256;row=row+1)
begin
col=col_row[row][s];
expanded_address=index_VN[row][col];
address_index=(col*2)+expanded_address;
AlphaSet[b][row]=doutA[address_index];
end
case(b)
QQ:state=`B_init2;
default:begin
a=a+1;
b=b+1;
end
endcase
end
`B_init2: begin
for(row=0;row<256;row=row+1) begin
col=col_row[row][s];
for(c = 0; c < (QQ+1); c=c+1)begin
						min_B[row][c] = max(AlphaSet[0][row],B[c][s+1][row]);

						for(b = 0; b < (QQ+1); b=b+1)begin
							mul_gf(H[row][col],b,mul_val);
                             add_gf(c,mul_val,a);

							max_B[row][c] = max(B[a][s + 1][row], AlphaSet[b][row]);
							min_B[row][c] = min(min_B[row][c], max_B[row][c]);

						end
						//B[c][s][row] = min_B[row][c];
						end
						end
						state=`B_init21;
						end
						`B_init21: begin
						for(row=0;row<256;row=row+1) begin
						for(c=0;c<(QQ+1);c=c+1) begin
						B[c][s][row] = min_B[row][c];
						end
						end
						
case(s)
1: begin
 s=0;
 state=`processing_state4;
end
0:begin
 state=`BETA1;
 a=0;
 end
endcase
end


`BETA1: begin
for(row=0;row<256;row=row+1)
begin
//for(a=0;a<4;a=a+1) begin
col=col_row[row][0];
expanded_address=index_CN[row][col];
address_index=(row*3);
addrBW[address_index]=a;
mul_gf(H[row][col],a,mul_val);
dinB[address_index]=B[mul_val][1][row];
weB[address_index]=1;
end
//end
for(row=0;row<256;row=row+1)
begin
//for(a=0;a<4;a=a+1) begin
col=col_row[row][2];
expanded_address=index_CN[row][col];
address_index=(row*3)+2;
addrBW[address_index]=a;
mul_gf(H[row][col],a,mul_val);
addrBW[address_index]=a;
dinB[address_index]=F[mul_val][1][row];
weB[address_index]=1;
end


for(row=0;row<256;row=row+1) begin
col=col_row[row][1];

                        mul_gf(H[row][col],a,mul_val);
						min_F[row][0] = max(F[mul_val][0][row], B[0][2][row]);

						for(b = 0; b < (QQ+1); b=b+1)begin
							mul_gf(H[row][col],a,mul_val);
                             add_gf(b,mul_val,c);
							max_F[row][0] = max(F[c][0][row],B[b][2][row]);

							min_F[row][0] = min(max_F[row][0], min_F[row][0]);

						end
						expanded_address=index_CN[row][col];
						address_index=(row*3)+1;
						addrBW[address_index]=a;
						dinB[address_index]=min_F[row][0];
						weB[address_index]=1;
end
case(a)
QQ:begin
state=`processing_state7;
c=0;
a=0;
end
default:
begin a=a+1;
end
endcase
end

 `processing_state7: begin
for(r=0;r<384;r=r+1)
begin
     
     row=row_col[1][r];//index1
     row_=row_col[0][r];//index0
     magicin=index_CN[row][r];//index1
     magic_=index_CN[row_][r];//index0
     m=magicin+(row*3);//index1
     p=magic_+(row_*3);//index0
     weB[m]=0;
     weB[p]=0;
     addrBR[m]=a;//index1
     addrBR[p]=a;//index0
     end       
 state=`s1;
 end
 `s1:begin
 state=`GammaFix;
 end
 
`GammaFix:begin
for(r=0;r<384;r=r+1)
begin
     row=row_col[1][r];//index1
     row_=row_col[0][r];//index0
     magicin=index_CN[row][r];//index1
     magic_=index_CN[row_][r];//index0
     m=magicin+(row*3);//index1
     p=magic_+(row_*3);//index0

tempa[a][r]=doutB[p]+Gamma[a][r];//indexv=0;
tempm[a][r]=doutB[m]+Gamma[a][r];//indexv=1
end
case(a)
QQ:begin
state=`s2;
a=0;
end
default:begin
a=a+1;
state=`processing_state7;
end
endcase
end     
          
`s2:begin
for(r=0;r<384;r=r+1)
begin
    minindex[0][r]=0;
    minindex[1][r]=2;
    minindex[2][r]=4;
    minindex[3][r]=6;
    for(a=0;a<2;a=a+1)
        begin
             if(tempa[a][r]<tempa[minindex[0][r]][r]) 
                minindex[0][r]=a;//index0
        end
    for(b=2;b<4;b=b+1)
        begin
             if(tempa[b][r]<tempa[minindex[1][r]][r]) 
                minindex[1][r]=b;//index0
        end    
        for(c=4;c<6;c=c+1)
        begin
             if(tempa[c][r]<tempa[minindex[2][r]][r]) 
                minindex[2][r]=c;//index0
        end    
         for(s=6;s<8;s=s+1)
        begin
             if(tempa[s][r]<tempa[minindex[3][r]][r]) 
                minindex[3][r]=s;//index0
        end    
        
     
             if(tempa[minindex[1][r]][r]<tempa[minindex[0][r]][r]) 
                minindex[0][r]=minindex[1][r];//index0
        //end    
       
             if(tempa[minindex[3][r]][r]<tempa[minindex[2][r]][r]) 
                minindex[2][r]=minindex[3][r];//index0
       // end    
  if(tempa[minindex[2][r]][r]<tempa[minindex[0][r]][r])
        minindex[0][r]=minindex[2][r];      
        end

for(t=0;t<384;t=t+1)
begin
 minindex_[0][t]=0;
    minindex_[1][t]=2;
    minindex_[2][t]=4;
    minindex_[3][t]=6;
    for(a=0;a<2;a=a+1)
        begin
             if(tempm[a][t]<tempm[minindex_[0][t]][t]) 
                minindex_[0][t]=a;//index1
        end
    for(b=2;b<4;b=b+1)
        begin
             if(tempm[b][t]<tempm[minindex_[1][t]][t]) 
                minindex_[1][t]=b;//index1
        end    
        for(c=4;c<6;c=c+1)
        begin
             if(tempm[c][t]<tempm[minindex_[2][t]][t]) 
                minindex_[2][t]=c;//index1
        end    
         for(s=6;s<8;s=s+1)
        begin
             if(tempm[s][t]<tempm[minindex_[3][t]][t]) 
                minindex_[3][t]=s;//index1
        end    
        
     
             if(tempm[minindex_[1][t]][t]<tempm[minindex_[0][t]][t]) 
                minindex_[0][t]=minindex_[1][t];//index1
        //end    
       
             if(tempm[minindex_[3][t]][t]<tempm[minindex_[2][t]][t]) 
                minindex_[2][t]=minindex_[3][t];//index1
       // end    
  if(tempm[minindex_[2][t]][t]<tempm[minindex_[0][t]][t])
        minindex_[0][t]=minindex_[2][t];      
       // end
        
        end
state=`FixAlpha;
a=0;
end

`FixAlpha:begin
 for(r=0;r<384;r=r+1)
     begin
     row=row_col[1][r];//index1
     magicin=index_VN[row][r];//1
     row_=row_col[0][r];//0
     magic_=index_VN[row_][r];//0
     p=magic_+(2*r);//0
     m=magicin+(2*r);//1
     addrAW[m]=a;//index1
     addrAW[p]=a;//index0
     weA[m]=1;
     weA[p]=1;
     dinA[p]=tempm[a][r]-tempm[minindex_[0][r]][r];//index0=index1
     dinA[m]=tempa[a][r]-tempa[minindex[0][r]][r];//index1=index0
     end
case(a)
QQ:begin
iter=iter-1;
    if(iter==0)
    state=`BETAOUT1;
    else
    state=`processing_statex;
 end   
default:begin
a=a+1;

end
endcase
end     


`BETAOUT1: begin
weB[0]=0;
addrBR[0]=0;
state=`BETAOUT2;

end
`BETAOUT2: begin
weB[0]=0;
addrBR[0]=1;
state=`BETAOUT;
address_index=0;
b=2;
//c=2;
address_index1=0;
end
		 
`BETAOUT: begin
beta=doutB[address_index];
addrBR[address_index1]=b;

case(b)
QQ: 
case(address_index1)
767: begin
state=`s39;
end
default: begin
b=0;
address_index1=address_index1+1;
end
endcase
1: begin
b=b+1;
address_index=address_index+1;
end
default: begin
b=b+1;
end
endcase
end

`s39: begin
end


endcase
end
end
endmodule